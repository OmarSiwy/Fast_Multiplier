//
// Bickerstaff Tree Compressor
// Algorithm: BICKERSTAFF
// Input Width: 64 bits
// Encoding: BOOTH
// Type: Signed
// Partial Products: 32
// Product Width: 128
// Reduction Stages: 8
//

module compressor_tree #(
    parameter PIPE = 0
)(
    input logic clk,
    input logic rst,
    input logic [64:0] pp [31:0],
    /* verilator lint_off ASCRANGE */
    input logic [31:0] cpl,
    /* verilator lint_on ASCRANGE */
    output logic [127:0] sum,
    output logic [127:0] carry
);
    localparam int COMPRESSOR_TREE_STAGES = PIPE ? 8 : 0;

    // FA and HA output wires
    logic fa_s0_c2_n0_s, fa_s0_c2_n0_c;
    logic fa_s0_c4_n1_s, fa_s0_c4_n1_c;
    logic fa_s0_c5_n2_s, fa_s0_c5_n2_c;
    logic fa_s0_c6_n3_s, fa_s0_c6_n3_c;
    logic fa_s0_c7_n4_s, fa_s0_c7_n4_c;
    logic fa_s0_c8_n5_s, fa_s0_c8_n5_c;
    logic fa_s0_c8_n6_s, fa_s0_c8_n6_c;
    logic fa_s0_c9_n7_s, fa_s0_c9_n7_c;
    logic fa_s0_c10_n8_s, fa_s0_c10_n8_c;
    logic fa_s0_c10_n9_s, fa_s0_c10_n9_c;
    logic fa_s0_c11_n10_s, fa_s0_c11_n10_c;
    logic fa_s0_c11_n11_s, fa_s0_c11_n11_c;
    logic fa_s0_c12_n12_s, fa_s0_c12_n12_c;
    logic fa_s0_c12_n13_s, fa_s0_c12_n13_c;
    logic fa_s0_c13_n14_s, fa_s0_c13_n14_c;
    logic fa_s0_c13_n15_s, fa_s0_c13_n15_c;
    logic fa_s0_c14_n16_s, fa_s0_c14_n16_c;
    logic fa_s0_c14_n17_s, fa_s0_c14_n17_c;
    logic fa_s0_c14_n18_s, fa_s0_c14_n18_c;
    logic fa_s0_c15_n19_s, fa_s0_c15_n19_c;
    logic fa_s0_c15_n20_s, fa_s0_c15_n20_c;
    logic fa_s0_c16_n21_s, fa_s0_c16_n21_c;
    logic fa_s0_c16_n22_s, fa_s0_c16_n22_c;
    logic fa_s0_c16_n23_s, fa_s0_c16_n23_c;
    logic fa_s0_c17_n24_s, fa_s0_c17_n24_c;
    logic fa_s0_c17_n25_s, fa_s0_c17_n25_c;
    logic fa_s0_c17_n26_s, fa_s0_c17_n26_c;
    logic fa_s0_c18_n27_s, fa_s0_c18_n27_c;
    logic fa_s0_c18_n28_s, fa_s0_c18_n28_c;
    logic fa_s0_c18_n29_s, fa_s0_c18_n29_c;
    logic fa_s0_c19_n30_s, fa_s0_c19_n30_c;
    logic fa_s0_c19_n31_s, fa_s0_c19_n31_c;
    logic fa_s0_c19_n32_s, fa_s0_c19_n32_c;
    logic fa_s0_c20_n33_s, fa_s0_c20_n33_c;
    logic fa_s0_c20_n34_s, fa_s0_c20_n34_c;
    logic fa_s0_c20_n35_s, fa_s0_c20_n35_c;
    logic fa_s0_c20_n36_s, fa_s0_c20_n36_c;
    logic fa_s0_c21_n37_s, fa_s0_c21_n37_c;
    logic fa_s0_c21_n38_s, fa_s0_c21_n38_c;
    logic fa_s0_c21_n39_s, fa_s0_c21_n39_c;
    logic fa_s0_c22_n40_s, fa_s0_c22_n40_c;
    logic fa_s0_c22_n41_s, fa_s0_c22_n41_c;
    logic fa_s0_c22_n42_s, fa_s0_c22_n42_c;
    logic fa_s0_c22_n43_s, fa_s0_c22_n43_c;
    logic fa_s0_c23_n44_s, fa_s0_c23_n44_c;
    logic fa_s0_c23_n45_s, fa_s0_c23_n45_c;
    logic fa_s0_c23_n46_s, fa_s0_c23_n46_c;
    logic fa_s0_c23_n47_s, fa_s0_c23_n47_c;
    logic fa_s0_c24_n48_s, fa_s0_c24_n48_c;
    logic fa_s0_c24_n49_s, fa_s0_c24_n49_c;
    logic fa_s0_c24_n50_s, fa_s0_c24_n50_c;
    logic fa_s0_c24_n51_s, fa_s0_c24_n51_c;
    logic fa_s0_c25_n52_s, fa_s0_c25_n52_c;
    logic fa_s0_c25_n53_s, fa_s0_c25_n53_c;
    logic fa_s0_c25_n54_s, fa_s0_c25_n54_c;
    logic fa_s0_c25_n55_s, fa_s0_c25_n55_c;
    logic fa_s0_c26_n56_s, fa_s0_c26_n56_c;
    logic fa_s0_c26_n57_s, fa_s0_c26_n57_c;
    logic fa_s0_c26_n58_s, fa_s0_c26_n58_c;
    logic fa_s0_c26_n59_s, fa_s0_c26_n59_c;
    logic fa_s0_c26_n60_s, fa_s0_c26_n60_c;
    logic fa_s0_c27_n61_s, fa_s0_c27_n61_c;
    logic fa_s0_c27_n62_s, fa_s0_c27_n62_c;
    logic fa_s0_c27_n63_s, fa_s0_c27_n63_c;
    logic fa_s0_c27_n64_s, fa_s0_c27_n64_c;
    logic fa_s0_c28_n65_s, fa_s0_c28_n65_c;
    logic fa_s0_c28_n66_s, fa_s0_c28_n66_c;
    logic fa_s0_c28_n67_s, fa_s0_c28_n67_c;
    logic fa_s0_c28_n68_s, fa_s0_c28_n68_c;
    logic fa_s0_c28_n69_s, fa_s0_c28_n69_c;
    logic fa_s0_c29_n70_s, fa_s0_c29_n70_c;
    logic fa_s0_c29_n71_s, fa_s0_c29_n71_c;
    logic fa_s0_c29_n72_s, fa_s0_c29_n72_c;
    logic fa_s0_c29_n73_s, fa_s0_c29_n73_c;
    logic fa_s0_c29_n74_s, fa_s0_c29_n74_c;
    logic fa_s0_c30_n75_s, fa_s0_c30_n75_c;
    logic fa_s0_c30_n76_s, fa_s0_c30_n76_c;
    logic fa_s0_c30_n77_s, fa_s0_c30_n77_c;
    logic fa_s0_c30_n78_s, fa_s0_c30_n78_c;
    logic fa_s0_c30_n79_s, fa_s0_c30_n79_c;
    logic fa_s0_c31_n80_s, fa_s0_c31_n80_c;
    logic fa_s0_c31_n81_s, fa_s0_c31_n81_c;
    logic fa_s0_c31_n82_s, fa_s0_c31_n82_c;
    logic fa_s0_c31_n83_s, fa_s0_c31_n83_c;
    logic fa_s0_c31_n84_s, fa_s0_c31_n84_c;
    logic fa_s0_c32_n85_s, fa_s0_c32_n85_c;
    logic fa_s0_c32_n86_s, fa_s0_c32_n86_c;
    logic fa_s0_c32_n87_s, fa_s0_c32_n87_c;
    logic fa_s0_c32_n88_s, fa_s0_c32_n88_c;
    logic fa_s0_c32_n89_s, fa_s0_c32_n89_c;
    logic fa_s0_c32_n90_s, fa_s0_c32_n90_c;
    logic fa_s0_c33_n91_s, fa_s0_c33_n91_c;
    logic fa_s0_c33_n92_s, fa_s0_c33_n92_c;
    logic fa_s0_c33_n93_s, fa_s0_c33_n93_c;
    logic fa_s0_c33_n94_s, fa_s0_c33_n94_c;
    logic fa_s0_c33_n95_s, fa_s0_c33_n95_c;
    logic fa_s0_c34_n96_s, fa_s0_c34_n96_c;
    logic fa_s0_c34_n97_s, fa_s0_c34_n97_c;
    logic fa_s0_c34_n98_s, fa_s0_c34_n98_c;
    logic fa_s0_c34_n99_s, fa_s0_c34_n99_c;
    logic fa_s0_c34_n100_s, fa_s0_c34_n100_c;
    logic fa_s0_c34_n101_s, fa_s0_c34_n101_c;
    logic fa_s0_c35_n102_s, fa_s0_c35_n102_c;
    logic fa_s0_c35_n103_s, fa_s0_c35_n103_c;
    logic fa_s0_c35_n104_s, fa_s0_c35_n104_c;
    logic fa_s0_c35_n105_s, fa_s0_c35_n105_c;
    logic fa_s0_c35_n106_s, fa_s0_c35_n106_c;
    logic fa_s0_c35_n107_s, fa_s0_c35_n107_c;
    logic fa_s0_c36_n108_s, fa_s0_c36_n108_c;
    logic fa_s0_c36_n109_s, fa_s0_c36_n109_c;
    logic fa_s0_c36_n110_s, fa_s0_c36_n110_c;
    logic fa_s0_c36_n111_s, fa_s0_c36_n111_c;
    logic fa_s0_c36_n112_s, fa_s0_c36_n112_c;
    logic fa_s0_c36_n113_s, fa_s0_c36_n113_c;
    logic fa_s0_c37_n114_s, fa_s0_c37_n114_c;
    logic fa_s0_c37_n115_s, fa_s0_c37_n115_c;
    logic fa_s0_c37_n116_s, fa_s0_c37_n116_c;
    logic fa_s0_c37_n117_s, fa_s0_c37_n117_c;
    logic fa_s0_c37_n118_s, fa_s0_c37_n118_c;
    logic fa_s0_c37_n119_s, fa_s0_c37_n119_c;
    logic fa_s0_c38_n120_s, fa_s0_c38_n120_c;
    logic fa_s0_c38_n121_s, fa_s0_c38_n121_c;
    logic fa_s0_c38_n122_s, fa_s0_c38_n122_c;
    logic fa_s0_c38_n123_s, fa_s0_c38_n123_c;
    logic fa_s0_c38_n124_s, fa_s0_c38_n124_c;
    logic fa_s0_c38_n125_s, fa_s0_c38_n125_c;
    logic fa_s0_c38_n126_s, fa_s0_c38_n126_c;
    logic fa_s0_c39_n127_s, fa_s0_c39_n127_c;
    logic fa_s0_c39_n128_s, fa_s0_c39_n128_c;
    logic fa_s0_c39_n129_s, fa_s0_c39_n129_c;
    logic fa_s0_c39_n130_s, fa_s0_c39_n130_c;
    logic fa_s0_c39_n131_s, fa_s0_c39_n131_c;
    logic fa_s0_c39_n132_s, fa_s0_c39_n132_c;
    logic fa_s0_c40_n133_s, fa_s0_c40_n133_c;
    logic fa_s0_c40_n134_s, fa_s0_c40_n134_c;
    logic fa_s0_c40_n135_s, fa_s0_c40_n135_c;
    logic fa_s0_c40_n136_s, fa_s0_c40_n136_c;
    logic fa_s0_c40_n137_s, fa_s0_c40_n137_c;
    logic fa_s0_c40_n138_s, fa_s0_c40_n138_c;
    logic fa_s0_c40_n139_s, fa_s0_c40_n139_c;
    logic fa_s0_c41_n140_s, fa_s0_c41_n140_c;
    logic fa_s0_c41_n141_s, fa_s0_c41_n141_c;
    logic fa_s0_c41_n142_s, fa_s0_c41_n142_c;
    logic fa_s0_c41_n143_s, fa_s0_c41_n143_c;
    logic fa_s0_c41_n144_s, fa_s0_c41_n144_c;
    logic fa_s0_c41_n145_s, fa_s0_c41_n145_c;
    logic fa_s0_c41_n146_s, fa_s0_c41_n146_c;
    logic fa_s0_c42_n147_s, fa_s0_c42_n147_c;
    logic fa_s0_c42_n148_s, fa_s0_c42_n148_c;
    logic fa_s0_c42_n149_s, fa_s0_c42_n149_c;
    logic fa_s0_c42_n150_s, fa_s0_c42_n150_c;
    logic fa_s0_c42_n151_s, fa_s0_c42_n151_c;
    logic fa_s0_c42_n152_s, fa_s0_c42_n152_c;
    logic fa_s0_c42_n153_s, fa_s0_c42_n153_c;
    logic fa_s0_c43_n154_s, fa_s0_c43_n154_c;
    logic fa_s0_c43_n155_s, fa_s0_c43_n155_c;
    logic fa_s0_c43_n156_s, fa_s0_c43_n156_c;
    logic fa_s0_c43_n157_s, fa_s0_c43_n157_c;
    logic fa_s0_c43_n158_s, fa_s0_c43_n158_c;
    logic fa_s0_c43_n159_s, fa_s0_c43_n159_c;
    logic fa_s0_c43_n160_s, fa_s0_c43_n160_c;
    logic fa_s0_c44_n161_s, fa_s0_c44_n161_c;
    logic fa_s0_c44_n162_s, fa_s0_c44_n162_c;
    logic fa_s0_c44_n163_s, fa_s0_c44_n163_c;
    logic fa_s0_c44_n164_s, fa_s0_c44_n164_c;
    logic fa_s0_c44_n165_s, fa_s0_c44_n165_c;
    logic fa_s0_c44_n166_s, fa_s0_c44_n166_c;
    logic fa_s0_c44_n167_s, fa_s0_c44_n167_c;
    logic fa_s0_c44_n168_s, fa_s0_c44_n168_c;
    logic fa_s0_c45_n169_s, fa_s0_c45_n169_c;
    logic fa_s0_c45_n170_s, fa_s0_c45_n170_c;
    logic fa_s0_c45_n171_s, fa_s0_c45_n171_c;
    logic fa_s0_c45_n172_s, fa_s0_c45_n172_c;
    logic fa_s0_c45_n173_s, fa_s0_c45_n173_c;
    logic fa_s0_c45_n174_s, fa_s0_c45_n174_c;
    logic fa_s0_c45_n175_s, fa_s0_c45_n175_c;
    logic fa_s0_c46_n176_s, fa_s0_c46_n176_c;
    logic fa_s0_c46_n177_s, fa_s0_c46_n177_c;
    logic fa_s0_c46_n178_s, fa_s0_c46_n178_c;
    logic fa_s0_c46_n179_s, fa_s0_c46_n179_c;
    logic fa_s0_c46_n180_s, fa_s0_c46_n180_c;
    logic fa_s0_c46_n181_s, fa_s0_c46_n181_c;
    logic fa_s0_c46_n182_s, fa_s0_c46_n182_c;
    logic fa_s0_c46_n183_s, fa_s0_c46_n183_c;
    logic fa_s0_c47_n184_s, fa_s0_c47_n184_c;
    logic fa_s0_c47_n185_s, fa_s0_c47_n185_c;
    logic fa_s0_c47_n186_s, fa_s0_c47_n186_c;
    logic fa_s0_c47_n187_s, fa_s0_c47_n187_c;
    logic fa_s0_c47_n188_s, fa_s0_c47_n188_c;
    logic fa_s0_c47_n189_s, fa_s0_c47_n189_c;
    logic fa_s0_c47_n190_s, fa_s0_c47_n190_c;
    logic fa_s0_c47_n191_s, fa_s0_c47_n191_c;
    logic fa_s0_c48_n192_s, fa_s0_c48_n192_c;
    logic fa_s0_c48_n193_s, fa_s0_c48_n193_c;
    logic fa_s0_c48_n194_s, fa_s0_c48_n194_c;
    logic fa_s0_c48_n195_s, fa_s0_c48_n195_c;
    logic fa_s0_c48_n196_s, fa_s0_c48_n196_c;
    logic fa_s0_c48_n197_s, fa_s0_c48_n197_c;
    logic fa_s0_c48_n198_s, fa_s0_c48_n198_c;
    logic fa_s0_c48_n199_s, fa_s0_c48_n199_c;
    logic fa_s0_c49_n200_s, fa_s0_c49_n200_c;
    logic fa_s0_c49_n201_s, fa_s0_c49_n201_c;
    logic fa_s0_c49_n202_s, fa_s0_c49_n202_c;
    logic fa_s0_c49_n203_s, fa_s0_c49_n203_c;
    logic fa_s0_c49_n204_s, fa_s0_c49_n204_c;
    logic fa_s0_c49_n205_s, fa_s0_c49_n205_c;
    logic fa_s0_c49_n206_s, fa_s0_c49_n206_c;
    logic fa_s0_c49_n207_s, fa_s0_c49_n207_c;
    logic fa_s0_c50_n208_s, fa_s0_c50_n208_c;
    logic fa_s0_c50_n209_s, fa_s0_c50_n209_c;
    logic fa_s0_c50_n210_s, fa_s0_c50_n210_c;
    logic fa_s0_c50_n211_s, fa_s0_c50_n211_c;
    logic fa_s0_c50_n212_s, fa_s0_c50_n212_c;
    logic fa_s0_c50_n213_s, fa_s0_c50_n213_c;
    logic fa_s0_c50_n214_s, fa_s0_c50_n214_c;
    logic fa_s0_c50_n215_s, fa_s0_c50_n215_c;
    logic fa_s0_c50_n216_s, fa_s0_c50_n216_c;
    logic fa_s0_c51_n217_s, fa_s0_c51_n217_c;
    logic fa_s0_c51_n218_s, fa_s0_c51_n218_c;
    logic fa_s0_c51_n219_s, fa_s0_c51_n219_c;
    logic fa_s0_c51_n220_s, fa_s0_c51_n220_c;
    logic fa_s0_c51_n221_s, fa_s0_c51_n221_c;
    logic fa_s0_c51_n222_s, fa_s0_c51_n222_c;
    logic fa_s0_c51_n223_s, fa_s0_c51_n223_c;
    logic fa_s0_c51_n224_s, fa_s0_c51_n224_c;
    logic fa_s0_c52_n225_s, fa_s0_c52_n225_c;
    logic fa_s0_c52_n226_s, fa_s0_c52_n226_c;
    logic fa_s0_c52_n227_s, fa_s0_c52_n227_c;
    logic fa_s0_c52_n228_s, fa_s0_c52_n228_c;
    logic fa_s0_c52_n229_s, fa_s0_c52_n229_c;
    logic fa_s0_c52_n230_s, fa_s0_c52_n230_c;
    logic fa_s0_c52_n231_s, fa_s0_c52_n231_c;
    logic fa_s0_c52_n232_s, fa_s0_c52_n232_c;
    logic fa_s0_c52_n233_s, fa_s0_c52_n233_c;
    logic fa_s0_c53_n234_s, fa_s0_c53_n234_c;
    logic fa_s0_c53_n235_s, fa_s0_c53_n235_c;
    logic fa_s0_c53_n236_s, fa_s0_c53_n236_c;
    logic fa_s0_c53_n237_s, fa_s0_c53_n237_c;
    logic fa_s0_c53_n238_s, fa_s0_c53_n238_c;
    logic fa_s0_c53_n239_s, fa_s0_c53_n239_c;
    logic fa_s0_c53_n240_s, fa_s0_c53_n240_c;
    logic fa_s0_c53_n241_s, fa_s0_c53_n241_c;
    logic fa_s0_c53_n242_s, fa_s0_c53_n242_c;
    logic fa_s0_c54_n243_s, fa_s0_c54_n243_c;
    logic fa_s0_c54_n244_s, fa_s0_c54_n244_c;
    logic fa_s0_c54_n245_s, fa_s0_c54_n245_c;
    logic fa_s0_c54_n246_s, fa_s0_c54_n246_c;
    logic fa_s0_c54_n247_s, fa_s0_c54_n247_c;
    logic fa_s0_c54_n248_s, fa_s0_c54_n248_c;
    logic fa_s0_c54_n249_s, fa_s0_c54_n249_c;
    logic fa_s0_c54_n250_s, fa_s0_c54_n250_c;
    logic fa_s0_c54_n251_s, fa_s0_c54_n251_c;
    logic fa_s0_c55_n252_s, fa_s0_c55_n252_c;
    logic fa_s0_c55_n253_s, fa_s0_c55_n253_c;
    logic fa_s0_c55_n254_s, fa_s0_c55_n254_c;
    logic fa_s0_c55_n255_s, fa_s0_c55_n255_c;
    logic fa_s0_c55_n256_s, fa_s0_c55_n256_c;
    logic fa_s0_c55_n257_s, fa_s0_c55_n257_c;
    logic fa_s0_c55_n258_s, fa_s0_c55_n258_c;
    logic fa_s0_c55_n259_s, fa_s0_c55_n259_c;
    logic fa_s0_c55_n260_s, fa_s0_c55_n260_c;
    logic fa_s0_c56_n261_s, fa_s0_c56_n261_c;
    logic fa_s0_c56_n262_s, fa_s0_c56_n262_c;
    logic fa_s0_c56_n263_s, fa_s0_c56_n263_c;
    logic fa_s0_c56_n264_s, fa_s0_c56_n264_c;
    logic fa_s0_c56_n265_s, fa_s0_c56_n265_c;
    logic fa_s0_c56_n266_s, fa_s0_c56_n266_c;
    logic fa_s0_c56_n267_s, fa_s0_c56_n267_c;
    logic fa_s0_c56_n268_s, fa_s0_c56_n268_c;
    logic fa_s0_c56_n269_s, fa_s0_c56_n269_c;
    logic fa_s0_c56_n270_s, fa_s0_c56_n270_c;
    logic fa_s0_c57_n271_s, fa_s0_c57_n271_c;
    logic fa_s0_c57_n272_s, fa_s0_c57_n272_c;
    logic fa_s0_c57_n273_s, fa_s0_c57_n273_c;
    logic fa_s0_c57_n274_s, fa_s0_c57_n274_c;
    logic fa_s0_c57_n275_s, fa_s0_c57_n275_c;
    logic fa_s0_c57_n276_s, fa_s0_c57_n276_c;
    logic fa_s0_c57_n277_s, fa_s0_c57_n277_c;
    logic fa_s0_c57_n278_s, fa_s0_c57_n278_c;
    logic fa_s0_c57_n279_s, fa_s0_c57_n279_c;
    logic fa_s0_c58_n280_s, fa_s0_c58_n280_c;
    logic fa_s0_c58_n281_s, fa_s0_c58_n281_c;
    logic fa_s0_c58_n282_s, fa_s0_c58_n282_c;
    logic fa_s0_c58_n283_s, fa_s0_c58_n283_c;
    logic fa_s0_c58_n284_s, fa_s0_c58_n284_c;
    logic fa_s0_c58_n285_s, fa_s0_c58_n285_c;
    logic fa_s0_c58_n286_s, fa_s0_c58_n286_c;
    logic fa_s0_c58_n287_s, fa_s0_c58_n287_c;
    logic fa_s0_c58_n288_s, fa_s0_c58_n288_c;
    logic fa_s0_c58_n289_s, fa_s0_c58_n289_c;
    logic fa_s0_c59_n290_s, fa_s0_c59_n290_c;
    logic fa_s0_c59_n291_s, fa_s0_c59_n291_c;
    logic fa_s0_c59_n292_s, fa_s0_c59_n292_c;
    logic fa_s0_c59_n293_s, fa_s0_c59_n293_c;
    logic fa_s0_c59_n294_s, fa_s0_c59_n294_c;
    logic fa_s0_c59_n295_s, fa_s0_c59_n295_c;
    logic fa_s0_c59_n296_s, fa_s0_c59_n296_c;
    logic fa_s0_c59_n297_s, fa_s0_c59_n297_c;
    logic fa_s0_c59_n298_s, fa_s0_c59_n298_c;
    logic fa_s0_c59_n299_s, fa_s0_c59_n299_c;
    logic fa_s0_c60_n300_s, fa_s0_c60_n300_c;
    logic fa_s0_c60_n301_s, fa_s0_c60_n301_c;
    logic fa_s0_c60_n302_s, fa_s0_c60_n302_c;
    logic fa_s0_c60_n303_s, fa_s0_c60_n303_c;
    logic fa_s0_c60_n304_s, fa_s0_c60_n304_c;
    logic fa_s0_c60_n305_s, fa_s0_c60_n305_c;
    logic fa_s0_c60_n306_s, fa_s0_c60_n306_c;
    logic fa_s0_c60_n307_s, fa_s0_c60_n307_c;
    logic fa_s0_c60_n308_s, fa_s0_c60_n308_c;
    logic fa_s0_c60_n309_s, fa_s0_c60_n309_c;
    logic fa_s0_c61_n310_s, fa_s0_c61_n310_c;
    logic fa_s0_c61_n311_s, fa_s0_c61_n311_c;
    logic fa_s0_c61_n312_s, fa_s0_c61_n312_c;
    logic fa_s0_c61_n313_s, fa_s0_c61_n313_c;
    logic fa_s0_c61_n314_s, fa_s0_c61_n314_c;
    logic fa_s0_c61_n315_s, fa_s0_c61_n315_c;
    logic fa_s0_c61_n316_s, fa_s0_c61_n316_c;
    logic fa_s0_c61_n317_s, fa_s0_c61_n317_c;
    logic fa_s0_c61_n318_s, fa_s0_c61_n318_c;
    logic fa_s0_c61_n319_s, fa_s0_c61_n319_c;
    logic fa_s0_c62_n320_s, fa_s0_c62_n320_c;
    logic fa_s0_c62_n321_s, fa_s0_c62_n321_c;
    logic fa_s0_c62_n322_s, fa_s0_c62_n322_c;
    logic fa_s0_c62_n323_s, fa_s0_c62_n323_c;
    logic fa_s0_c62_n324_s, fa_s0_c62_n324_c;
    logic fa_s0_c62_n325_s, fa_s0_c62_n325_c;
    logic fa_s0_c62_n326_s, fa_s0_c62_n326_c;
    logic fa_s0_c62_n327_s, fa_s0_c62_n327_c;
    logic fa_s0_c62_n328_s, fa_s0_c62_n328_c;
    logic fa_s0_c62_n329_s, fa_s0_c62_n329_c;
    logic fa_s0_c62_n330_s, fa_s0_c62_n330_c;
    logic fa_s0_c63_n331_s, fa_s0_c63_n331_c;
    logic fa_s0_c63_n332_s, fa_s0_c63_n332_c;
    logic fa_s0_c63_n333_s, fa_s0_c63_n333_c;
    logic fa_s0_c63_n334_s, fa_s0_c63_n334_c;
    logic fa_s0_c63_n335_s, fa_s0_c63_n335_c;
    logic fa_s0_c63_n336_s, fa_s0_c63_n336_c;
    logic fa_s0_c63_n337_s, fa_s0_c63_n337_c;
    logic fa_s0_c63_n338_s, fa_s0_c63_n338_c;
    logic fa_s0_c63_n339_s, fa_s0_c63_n339_c;
    logic fa_s0_c63_n340_s, fa_s0_c63_n340_c;
    logic fa_s0_c64_n341_s, fa_s0_c64_n341_c;
    logic fa_s0_c64_n342_s, fa_s0_c64_n342_c;
    logic fa_s0_c64_n343_s, fa_s0_c64_n343_c;
    logic fa_s0_c64_n344_s, fa_s0_c64_n344_c;
    logic fa_s0_c64_n345_s, fa_s0_c64_n345_c;
    logic fa_s0_c64_n346_s, fa_s0_c64_n346_c;
    logic fa_s0_c64_n347_s, fa_s0_c64_n347_c;
    logic fa_s0_c64_n348_s, fa_s0_c64_n348_c;
    logic fa_s0_c64_n349_s, fa_s0_c64_n349_c;
    logic fa_s0_c64_n350_s, fa_s0_c64_n350_c;
    logic fa_s0_c64_n351_s, fa_s0_c64_n351_c;
    logic fa_s0_c65_n352_s, fa_s0_c65_n352_c;
    logic fa_s0_c65_n353_s, fa_s0_c65_n353_c;
    logic fa_s0_c65_n354_s, fa_s0_c65_n354_c;
    logic fa_s0_c65_n355_s, fa_s0_c65_n355_c;
    logic fa_s0_c65_n356_s, fa_s0_c65_n356_c;
    logic fa_s0_c65_n357_s, fa_s0_c65_n357_c;
    logic fa_s0_c65_n358_s, fa_s0_c65_n358_c;
    logic fa_s0_c65_n359_s, fa_s0_c65_n359_c;
    logic fa_s0_c65_n360_s, fa_s0_c65_n360_c;
    logic fa_s0_c65_n361_s, fa_s0_c65_n361_c;
    logic fa_s0_c66_n362_s, fa_s0_c66_n362_c;
    logic fa_s0_c66_n363_s, fa_s0_c66_n363_c;
    logic fa_s0_c66_n364_s, fa_s0_c66_n364_c;
    logic fa_s0_c66_n365_s, fa_s0_c66_n365_c;
    logic fa_s0_c66_n366_s, fa_s0_c66_n366_c;
    logic fa_s0_c66_n367_s, fa_s0_c66_n367_c;
    logic fa_s0_c66_n368_s, fa_s0_c66_n368_c;
    logic fa_s0_c66_n369_s, fa_s0_c66_n369_c;
    logic fa_s0_c66_n370_s, fa_s0_c66_n370_c;
    logic fa_s0_c66_n371_s, fa_s0_c66_n371_c;
    logic fa_s0_c66_n372_s, fa_s0_c66_n372_c;
    logic fa_s0_c67_n373_s, fa_s0_c67_n373_c;
    logic fa_s0_c67_n374_s, fa_s0_c67_n374_c;
    logic fa_s0_c67_n375_s, fa_s0_c67_n375_c;
    logic fa_s0_c67_n376_s, fa_s0_c67_n376_c;
    logic fa_s0_c67_n377_s, fa_s0_c67_n377_c;
    logic fa_s0_c67_n378_s, fa_s0_c67_n378_c;
    logic fa_s0_c67_n379_s, fa_s0_c67_n379_c;
    logic fa_s0_c67_n380_s, fa_s0_c67_n380_c;
    logic fa_s0_c67_n381_s, fa_s0_c67_n381_c;
    logic fa_s0_c67_n382_s, fa_s0_c67_n382_c;
    logic fa_s0_c68_n383_s, fa_s0_c68_n383_c;
    logic fa_s0_c68_n384_s, fa_s0_c68_n384_c;
    logic fa_s0_c68_n385_s, fa_s0_c68_n385_c;
    logic fa_s0_c68_n386_s, fa_s0_c68_n386_c;
    logic fa_s0_c68_n387_s, fa_s0_c68_n387_c;
    logic fa_s0_c68_n388_s, fa_s0_c68_n388_c;
    logic fa_s0_c68_n389_s, fa_s0_c68_n389_c;
    logic fa_s0_c68_n390_s, fa_s0_c68_n390_c;
    logic fa_s0_c68_n391_s, fa_s0_c68_n391_c;
    logic fa_s0_c68_n392_s, fa_s0_c68_n392_c;
    logic fa_s0_c68_n393_s, fa_s0_c68_n393_c;
    logic fa_s0_c69_n394_s, fa_s0_c69_n394_c;
    logic fa_s0_c69_n395_s, fa_s0_c69_n395_c;
    logic fa_s0_c69_n396_s, fa_s0_c69_n396_c;
    logic fa_s0_c69_n397_s, fa_s0_c69_n397_c;
    logic fa_s0_c69_n398_s, fa_s0_c69_n398_c;
    logic fa_s0_c69_n399_s, fa_s0_c69_n399_c;
    logic fa_s0_c69_n400_s, fa_s0_c69_n400_c;
    logic fa_s0_c69_n401_s, fa_s0_c69_n401_c;
    logic fa_s0_c69_n402_s, fa_s0_c69_n402_c;
    logic fa_s0_c69_n403_s, fa_s0_c69_n403_c;
    logic fa_s0_c70_n404_s, fa_s0_c70_n404_c;
    logic fa_s0_c70_n405_s, fa_s0_c70_n405_c;
    logic fa_s0_c70_n406_s, fa_s0_c70_n406_c;
    logic fa_s0_c70_n407_s, fa_s0_c70_n407_c;
    logic fa_s0_c70_n408_s, fa_s0_c70_n408_c;
    logic fa_s0_c70_n409_s, fa_s0_c70_n409_c;
    logic fa_s0_c70_n410_s, fa_s0_c70_n410_c;
    logic fa_s0_c70_n411_s, fa_s0_c70_n411_c;
    logic fa_s0_c70_n412_s, fa_s0_c70_n412_c;
    logic fa_s0_c70_n413_s, fa_s0_c70_n413_c;
    logic fa_s0_c70_n414_s, fa_s0_c70_n414_c;
    logic fa_s0_c71_n415_s, fa_s0_c71_n415_c;
    logic fa_s0_c71_n416_s, fa_s0_c71_n416_c;
    logic fa_s0_c71_n417_s, fa_s0_c71_n417_c;
    logic fa_s0_c71_n418_s, fa_s0_c71_n418_c;
    logic fa_s0_c71_n419_s, fa_s0_c71_n419_c;
    logic fa_s0_c71_n420_s, fa_s0_c71_n420_c;
    logic fa_s0_c71_n421_s, fa_s0_c71_n421_c;
    logic fa_s0_c71_n422_s, fa_s0_c71_n422_c;
    logic fa_s0_c71_n423_s, fa_s0_c71_n423_c;
    logic fa_s0_c71_n424_s, fa_s0_c71_n424_c;
    logic fa_s0_c72_n425_s, fa_s0_c72_n425_c;
    logic fa_s0_c72_n426_s, fa_s0_c72_n426_c;
    logic fa_s0_c72_n427_s, fa_s0_c72_n427_c;
    logic fa_s0_c72_n428_s, fa_s0_c72_n428_c;
    logic fa_s0_c72_n429_s, fa_s0_c72_n429_c;
    logic fa_s0_c72_n430_s, fa_s0_c72_n430_c;
    logic fa_s0_c72_n431_s, fa_s0_c72_n431_c;
    logic fa_s0_c72_n432_s, fa_s0_c72_n432_c;
    logic fa_s0_c72_n433_s, fa_s0_c72_n433_c;
    logic fa_s0_c72_n434_s, fa_s0_c72_n434_c;
    logic fa_s0_c72_n435_s, fa_s0_c72_n435_c;
    logic fa_s0_c73_n436_s, fa_s0_c73_n436_c;
    logic fa_s0_c73_n437_s, fa_s0_c73_n437_c;
    logic fa_s0_c73_n438_s, fa_s0_c73_n438_c;
    logic fa_s0_c73_n439_s, fa_s0_c73_n439_c;
    logic fa_s0_c73_n440_s, fa_s0_c73_n440_c;
    logic fa_s0_c73_n441_s, fa_s0_c73_n441_c;
    logic fa_s0_c73_n442_s, fa_s0_c73_n442_c;
    logic fa_s0_c73_n443_s, fa_s0_c73_n443_c;
    logic fa_s0_c73_n444_s, fa_s0_c73_n444_c;
    logic fa_s0_c73_n445_s, fa_s0_c73_n445_c;
    logic fa_s0_c74_n446_s, fa_s0_c74_n446_c;
    logic fa_s0_c74_n447_s, fa_s0_c74_n447_c;
    logic fa_s0_c74_n448_s, fa_s0_c74_n448_c;
    logic fa_s0_c74_n449_s, fa_s0_c74_n449_c;
    logic fa_s0_c74_n450_s, fa_s0_c74_n450_c;
    logic fa_s0_c74_n451_s, fa_s0_c74_n451_c;
    logic fa_s0_c74_n452_s, fa_s0_c74_n452_c;
    logic fa_s0_c74_n453_s, fa_s0_c74_n453_c;
    logic fa_s0_c74_n454_s, fa_s0_c74_n454_c;
    logic fa_s0_c74_n455_s, fa_s0_c74_n455_c;
    logic fa_s0_c74_n456_s, fa_s0_c74_n456_c;
    logic fa_s0_c75_n457_s, fa_s0_c75_n457_c;
    logic fa_s0_c75_n458_s, fa_s0_c75_n458_c;
    logic fa_s0_c75_n459_s, fa_s0_c75_n459_c;
    logic fa_s0_c75_n460_s, fa_s0_c75_n460_c;
    logic fa_s0_c75_n461_s, fa_s0_c75_n461_c;
    logic fa_s0_c75_n462_s, fa_s0_c75_n462_c;
    logic fa_s0_c75_n463_s, fa_s0_c75_n463_c;
    logic fa_s0_c75_n464_s, fa_s0_c75_n464_c;
    logic fa_s0_c75_n465_s, fa_s0_c75_n465_c;
    logic fa_s0_c75_n466_s, fa_s0_c75_n466_c;
    logic fa_s0_c76_n467_s, fa_s0_c76_n467_c;
    logic fa_s0_c76_n468_s, fa_s0_c76_n468_c;
    logic fa_s0_c76_n469_s, fa_s0_c76_n469_c;
    logic fa_s0_c76_n470_s, fa_s0_c76_n470_c;
    logic fa_s0_c76_n471_s, fa_s0_c76_n471_c;
    logic fa_s0_c76_n472_s, fa_s0_c76_n472_c;
    logic fa_s0_c76_n473_s, fa_s0_c76_n473_c;
    logic fa_s0_c76_n474_s, fa_s0_c76_n474_c;
    logic fa_s0_c76_n475_s, fa_s0_c76_n475_c;
    logic fa_s0_c76_n476_s, fa_s0_c76_n476_c;
    logic fa_s0_c76_n477_s, fa_s0_c76_n477_c;
    logic fa_s0_c77_n478_s, fa_s0_c77_n478_c;
    logic fa_s0_c77_n479_s, fa_s0_c77_n479_c;
    logic fa_s0_c77_n480_s, fa_s0_c77_n480_c;
    logic fa_s0_c77_n481_s, fa_s0_c77_n481_c;
    logic fa_s0_c77_n482_s, fa_s0_c77_n482_c;
    logic fa_s0_c77_n483_s, fa_s0_c77_n483_c;
    logic fa_s0_c77_n484_s, fa_s0_c77_n484_c;
    logic fa_s0_c77_n485_s, fa_s0_c77_n485_c;
    logic fa_s0_c77_n486_s, fa_s0_c77_n486_c;
    logic fa_s0_c77_n487_s, fa_s0_c77_n487_c;
    logic fa_s0_c78_n488_s, fa_s0_c78_n488_c;
    logic fa_s0_c78_n489_s, fa_s0_c78_n489_c;
    logic fa_s0_c78_n490_s, fa_s0_c78_n490_c;
    logic fa_s0_c78_n491_s, fa_s0_c78_n491_c;
    logic fa_s0_c78_n492_s, fa_s0_c78_n492_c;
    logic fa_s0_c78_n493_s, fa_s0_c78_n493_c;
    logic fa_s0_c78_n494_s, fa_s0_c78_n494_c;
    logic fa_s0_c78_n495_s, fa_s0_c78_n495_c;
    logic fa_s0_c78_n496_s, fa_s0_c78_n496_c;
    logic fa_s0_c78_n497_s, fa_s0_c78_n497_c;
    logic fa_s0_c78_n498_s, fa_s0_c78_n498_c;
    logic fa_s0_c79_n499_s, fa_s0_c79_n499_c;
    logic fa_s0_c79_n500_s, fa_s0_c79_n500_c;
    logic fa_s0_c79_n501_s, fa_s0_c79_n501_c;
    logic fa_s0_c79_n502_s, fa_s0_c79_n502_c;
    logic fa_s0_c79_n503_s, fa_s0_c79_n503_c;
    logic fa_s0_c79_n504_s, fa_s0_c79_n504_c;
    logic fa_s0_c79_n505_s, fa_s0_c79_n505_c;
    logic fa_s0_c79_n506_s, fa_s0_c79_n506_c;
    logic fa_s0_c79_n507_s, fa_s0_c79_n507_c;
    logic fa_s0_c79_n508_s, fa_s0_c79_n508_c;
    logic fa_s0_c80_n509_s, fa_s0_c80_n509_c;
    logic fa_s0_c80_n510_s, fa_s0_c80_n510_c;
    logic fa_s0_c80_n511_s, fa_s0_c80_n511_c;
    logic fa_s0_c80_n512_s, fa_s0_c80_n512_c;
    logic fa_s0_c80_n513_s, fa_s0_c80_n513_c;
    logic fa_s0_c80_n514_s, fa_s0_c80_n514_c;
    logic fa_s0_c80_n515_s, fa_s0_c80_n515_c;
    logic fa_s0_c80_n516_s, fa_s0_c80_n516_c;
    logic fa_s0_c80_n517_s, fa_s0_c80_n517_c;
    logic fa_s0_c80_n518_s, fa_s0_c80_n518_c;
    logic fa_s0_c80_n519_s, fa_s0_c80_n519_c;
    logic fa_s0_c81_n520_s, fa_s0_c81_n520_c;
    logic fa_s0_c81_n521_s, fa_s0_c81_n521_c;
    logic fa_s0_c81_n522_s, fa_s0_c81_n522_c;
    logic fa_s0_c81_n523_s, fa_s0_c81_n523_c;
    logic fa_s0_c81_n524_s, fa_s0_c81_n524_c;
    logic fa_s0_c81_n525_s, fa_s0_c81_n525_c;
    logic fa_s0_c81_n526_s, fa_s0_c81_n526_c;
    logic fa_s0_c81_n527_s, fa_s0_c81_n527_c;
    logic fa_s0_c81_n528_s, fa_s0_c81_n528_c;
    logic fa_s0_c81_n529_s, fa_s0_c81_n529_c;
    logic fa_s0_c82_n530_s, fa_s0_c82_n530_c;
    logic fa_s0_c82_n531_s, fa_s0_c82_n531_c;
    logic fa_s0_c82_n532_s, fa_s0_c82_n532_c;
    logic fa_s0_c82_n533_s, fa_s0_c82_n533_c;
    logic fa_s0_c82_n534_s, fa_s0_c82_n534_c;
    logic fa_s0_c82_n535_s, fa_s0_c82_n535_c;
    logic fa_s0_c82_n536_s, fa_s0_c82_n536_c;
    logic fa_s0_c82_n537_s, fa_s0_c82_n537_c;
    logic fa_s0_c82_n538_s, fa_s0_c82_n538_c;
    logic fa_s0_c82_n539_s, fa_s0_c82_n539_c;
    logic fa_s0_c82_n540_s, fa_s0_c82_n540_c;
    logic fa_s0_c83_n541_s, fa_s0_c83_n541_c;
    logic fa_s0_c83_n542_s, fa_s0_c83_n542_c;
    logic fa_s0_c83_n543_s, fa_s0_c83_n543_c;
    logic fa_s0_c83_n544_s, fa_s0_c83_n544_c;
    logic fa_s0_c83_n545_s, fa_s0_c83_n545_c;
    logic fa_s0_c83_n546_s, fa_s0_c83_n546_c;
    logic fa_s0_c83_n547_s, fa_s0_c83_n547_c;
    logic fa_s0_c83_n548_s, fa_s0_c83_n548_c;
    logic fa_s0_c83_n549_s, fa_s0_c83_n549_c;
    logic fa_s0_c83_n550_s, fa_s0_c83_n550_c;
    logic fa_s0_c84_n551_s, fa_s0_c84_n551_c;
    logic fa_s0_c84_n552_s, fa_s0_c84_n552_c;
    logic fa_s0_c84_n553_s, fa_s0_c84_n553_c;
    logic fa_s0_c84_n554_s, fa_s0_c84_n554_c;
    logic fa_s0_c84_n555_s, fa_s0_c84_n555_c;
    logic fa_s0_c84_n556_s, fa_s0_c84_n556_c;
    logic fa_s0_c84_n557_s, fa_s0_c84_n557_c;
    logic fa_s0_c84_n558_s, fa_s0_c84_n558_c;
    logic fa_s0_c84_n559_s, fa_s0_c84_n559_c;
    logic fa_s0_c84_n560_s, fa_s0_c84_n560_c;
    logic fa_s0_c84_n561_s, fa_s0_c84_n561_c;
    logic fa_s0_c85_n562_s, fa_s0_c85_n562_c;
    logic fa_s0_c85_n563_s, fa_s0_c85_n563_c;
    logic fa_s0_c85_n564_s, fa_s0_c85_n564_c;
    logic fa_s0_c85_n565_s, fa_s0_c85_n565_c;
    logic fa_s0_c85_n566_s, fa_s0_c85_n566_c;
    logic fa_s0_c85_n567_s, fa_s0_c85_n567_c;
    logic fa_s0_c85_n568_s, fa_s0_c85_n568_c;
    logic fa_s0_c85_n569_s, fa_s0_c85_n569_c;
    logic fa_s0_c85_n570_s, fa_s0_c85_n570_c;
    logic fa_s0_c85_n571_s, fa_s0_c85_n571_c;
    logic fa_s0_c86_n572_s, fa_s0_c86_n572_c;
    logic fa_s0_c86_n573_s, fa_s0_c86_n573_c;
    logic fa_s0_c86_n574_s, fa_s0_c86_n574_c;
    logic fa_s0_c86_n575_s, fa_s0_c86_n575_c;
    logic fa_s0_c86_n576_s, fa_s0_c86_n576_c;
    logic fa_s0_c86_n577_s, fa_s0_c86_n577_c;
    logic fa_s0_c86_n578_s, fa_s0_c86_n578_c;
    logic fa_s0_c86_n579_s, fa_s0_c86_n579_c;
    logic fa_s0_c86_n580_s, fa_s0_c86_n580_c;
    logic fa_s0_c86_n581_s, fa_s0_c86_n581_c;
    logic fa_s0_c86_n582_s, fa_s0_c86_n582_c;
    logic fa_s0_c87_n583_s, fa_s0_c87_n583_c;
    logic fa_s0_c87_n584_s, fa_s0_c87_n584_c;
    logic fa_s0_c87_n585_s, fa_s0_c87_n585_c;
    logic fa_s0_c87_n586_s, fa_s0_c87_n586_c;
    logic fa_s0_c87_n587_s, fa_s0_c87_n587_c;
    logic fa_s0_c87_n588_s, fa_s0_c87_n588_c;
    logic fa_s0_c87_n589_s, fa_s0_c87_n589_c;
    logic fa_s0_c87_n590_s, fa_s0_c87_n590_c;
    logic fa_s0_c87_n591_s, fa_s0_c87_n591_c;
    logic fa_s0_c87_n592_s, fa_s0_c87_n592_c;
    logic fa_s0_c88_n593_s, fa_s0_c88_n593_c;
    logic fa_s0_c88_n594_s, fa_s0_c88_n594_c;
    logic fa_s0_c88_n595_s, fa_s0_c88_n595_c;
    logic fa_s0_c88_n596_s, fa_s0_c88_n596_c;
    logic fa_s0_c88_n597_s, fa_s0_c88_n597_c;
    logic fa_s0_c88_n598_s, fa_s0_c88_n598_c;
    logic fa_s0_c88_n599_s, fa_s0_c88_n599_c;
    logic fa_s0_c88_n600_s, fa_s0_c88_n600_c;
    logic fa_s0_c88_n601_s, fa_s0_c88_n601_c;
    logic fa_s0_c88_n602_s, fa_s0_c88_n602_c;
    logic fa_s0_c88_n603_s, fa_s0_c88_n603_c;
    logic fa_s0_c89_n604_s, fa_s0_c89_n604_c;
    logic fa_s0_c89_n605_s, fa_s0_c89_n605_c;
    logic fa_s0_c89_n606_s, fa_s0_c89_n606_c;
    logic fa_s0_c89_n607_s, fa_s0_c89_n607_c;
    logic fa_s0_c89_n608_s, fa_s0_c89_n608_c;
    logic fa_s0_c89_n609_s, fa_s0_c89_n609_c;
    logic fa_s0_c89_n610_s, fa_s0_c89_n610_c;
    logic fa_s0_c89_n611_s, fa_s0_c89_n611_c;
    logic fa_s0_c89_n612_s, fa_s0_c89_n612_c;
    logic fa_s0_c89_n613_s, fa_s0_c89_n613_c;
    logic fa_s0_c90_n614_s, fa_s0_c90_n614_c;
    logic fa_s0_c90_n615_s, fa_s0_c90_n615_c;
    logic fa_s0_c90_n616_s, fa_s0_c90_n616_c;
    logic fa_s0_c90_n617_s, fa_s0_c90_n617_c;
    logic fa_s0_c90_n618_s, fa_s0_c90_n618_c;
    logic fa_s0_c90_n619_s, fa_s0_c90_n619_c;
    logic fa_s0_c90_n620_s, fa_s0_c90_n620_c;
    logic fa_s0_c90_n621_s, fa_s0_c90_n621_c;
    logic fa_s0_c90_n622_s, fa_s0_c90_n622_c;
    logic fa_s0_c90_n623_s, fa_s0_c90_n623_c;
    logic fa_s0_c90_n624_s, fa_s0_c90_n624_c;
    logic fa_s0_c91_n625_s, fa_s0_c91_n625_c;
    logic fa_s0_c91_n626_s, fa_s0_c91_n626_c;
    logic fa_s0_c91_n627_s, fa_s0_c91_n627_c;
    logic fa_s0_c91_n628_s, fa_s0_c91_n628_c;
    logic fa_s0_c91_n629_s, fa_s0_c91_n629_c;
    logic fa_s0_c91_n630_s, fa_s0_c91_n630_c;
    logic fa_s0_c91_n631_s, fa_s0_c91_n631_c;
    logic fa_s0_c91_n632_s, fa_s0_c91_n632_c;
    logic fa_s0_c91_n633_s, fa_s0_c91_n633_c;
    logic fa_s0_c91_n634_s, fa_s0_c91_n634_c;
    logic fa_s0_c92_n635_s, fa_s0_c92_n635_c;
    logic fa_s0_c92_n636_s, fa_s0_c92_n636_c;
    logic fa_s0_c92_n637_s, fa_s0_c92_n637_c;
    logic fa_s0_c92_n638_s, fa_s0_c92_n638_c;
    logic fa_s0_c92_n639_s, fa_s0_c92_n639_c;
    logic fa_s0_c92_n640_s, fa_s0_c92_n640_c;
    logic fa_s0_c92_n641_s, fa_s0_c92_n641_c;
    logic fa_s0_c92_n642_s, fa_s0_c92_n642_c;
    logic fa_s0_c92_n643_s, fa_s0_c92_n643_c;
    logic fa_s0_c92_n644_s, fa_s0_c92_n644_c;
    logic fa_s0_c92_n645_s, fa_s0_c92_n645_c;
    logic fa_s0_c93_n646_s, fa_s0_c93_n646_c;
    logic fa_s0_c93_n647_s, fa_s0_c93_n647_c;
    logic fa_s0_c93_n648_s, fa_s0_c93_n648_c;
    logic fa_s0_c93_n649_s, fa_s0_c93_n649_c;
    logic fa_s0_c93_n650_s, fa_s0_c93_n650_c;
    logic fa_s0_c93_n651_s, fa_s0_c93_n651_c;
    logic fa_s0_c93_n652_s, fa_s0_c93_n652_c;
    logic fa_s0_c93_n653_s, fa_s0_c93_n653_c;
    logic fa_s0_c93_n654_s, fa_s0_c93_n654_c;
    logic fa_s0_c93_n655_s, fa_s0_c93_n655_c;
    logic fa_s0_c94_n656_s, fa_s0_c94_n656_c;
    logic fa_s0_c94_n657_s, fa_s0_c94_n657_c;
    logic fa_s0_c94_n658_s, fa_s0_c94_n658_c;
    logic fa_s0_c94_n659_s, fa_s0_c94_n659_c;
    logic fa_s0_c94_n660_s, fa_s0_c94_n660_c;
    logic fa_s0_c94_n661_s, fa_s0_c94_n661_c;
    logic fa_s0_c94_n662_s, fa_s0_c94_n662_c;
    logic fa_s0_c94_n663_s, fa_s0_c94_n663_c;
    logic fa_s0_c94_n664_s, fa_s0_c94_n664_c;
    logic fa_s0_c94_n665_s, fa_s0_c94_n665_c;
    logic fa_s0_c94_n666_s, fa_s0_c94_n666_c;
    logic fa_s0_c95_n667_s, fa_s0_c95_n667_c;
    logic fa_s0_c95_n668_s, fa_s0_c95_n668_c;
    logic fa_s0_c95_n669_s, fa_s0_c95_n669_c;
    logic fa_s0_c95_n670_s, fa_s0_c95_n670_c;
    logic fa_s0_c95_n671_s, fa_s0_c95_n671_c;
    logic fa_s0_c95_n672_s, fa_s0_c95_n672_c;
    logic fa_s0_c95_n673_s, fa_s0_c95_n673_c;
    logic fa_s0_c95_n674_s, fa_s0_c95_n674_c;
    logic fa_s0_c95_n675_s, fa_s0_c95_n675_c;
    logic fa_s0_c95_n676_s, fa_s0_c95_n676_c;
    logic fa_s0_c96_n677_s, fa_s0_c96_n677_c;
    logic fa_s0_c96_n678_s, fa_s0_c96_n678_c;
    logic fa_s0_c96_n679_s, fa_s0_c96_n679_c;
    logic fa_s0_c96_n680_s, fa_s0_c96_n680_c;
    logic fa_s0_c96_n681_s, fa_s0_c96_n681_c;
    logic fa_s0_c96_n682_s, fa_s0_c96_n682_c;
    logic fa_s0_c96_n683_s, fa_s0_c96_n683_c;
    logic fa_s0_c96_n684_s, fa_s0_c96_n684_c;
    logic fa_s0_c96_n685_s, fa_s0_c96_n685_c;
    logic fa_s0_c96_n686_s, fa_s0_c96_n686_c;
    logic fa_s0_c96_n687_s, fa_s0_c96_n687_c;
    logic fa_s0_c97_n688_s, fa_s0_c97_n688_c;
    logic fa_s0_c97_n689_s, fa_s0_c97_n689_c;
    logic fa_s0_c97_n690_s, fa_s0_c97_n690_c;
    logic fa_s0_c97_n691_s, fa_s0_c97_n691_c;
    logic fa_s0_c97_n692_s, fa_s0_c97_n692_c;
    logic fa_s0_c97_n693_s, fa_s0_c97_n693_c;
    logic fa_s0_c97_n694_s, fa_s0_c97_n694_c;
    logic fa_s0_c97_n695_s, fa_s0_c97_n695_c;
    logic fa_s0_c97_n696_s, fa_s0_c97_n696_c;
    logic fa_s0_c97_n697_s, fa_s0_c97_n697_c;
    logic fa_s0_c98_n698_s, fa_s0_c98_n698_c;
    logic fa_s0_c98_n699_s, fa_s0_c98_n699_c;
    logic fa_s0_c98_n700_s, fa_s0_c98_n700_c;
    logic fa_s0_c98_n701_s, fa_s0_c98_n701_c;
    logic fa_s0_c98_n702_s, fa_s0_c98_n702_c;
    logic fa_s0_c98_n703_s, fa_s0_c98_n703_c;
    logic fa_s0_c98_n704_s, fa_s0_c98_n704_c;
    logic fa_s0_c98_n705_s, fa_s0_c98_n705_c;
    logic fa_s0_c98_n706_s, fa_s0_c98_n706_c;
    logic fa_s0_c98_n707_s, fa_s0_c98_n707_c;
    logic fa_s0_c98_n708_s, fa_s0_c98_n708_c;
    logic fa_s0_c99_n709_s, fa_s0_c99_n709_c;
    logic fa_s0_c99_n710_s, fa_s0_c99_n710_c;
    logic fa_s0_c99_n711_s, fa_s0_c99_n711_c;
    logic fa_s0_c99_n712_s, fa_s0_c99_n712_c;
    logic fa_s0_c99_n713_s, fa_s0_c99_n713_c;
    logic fa_s0_c99_n714_s, fa_s0_c99_n714_c;
    logic fa_s0_c99_n715_s, fa_s0_c99_n715_c;
    logic fa_s0_c99_n716_s, fa_s0_c99_n716_c;
    logic fa_s0_c99_n717_s, fa_s0_c99_n717_c;
    logic fa_s0_c99_n718_s, fa_s0_c99_n718_c;
    logic fa_s0_c100_n719_s, fa_s0_c100_n719_c;
    logic fa_s0_c100_n720_s, fa_s0_c100_n720_c;
    logic fa_s0_c100_n721_s, fa_s0_c100_n721_c;
    logic fa_s0_c100_n722_s, fa_s0_c100_n722_c;
    logic fa_s0_c100_n723_s, fa_s0_c100_n723_c;
    logic fa_s0_c100_n724_s, fa_s0_c100_n724_c;
    logic fa_s0_c100_n725_s, fa_s0_c100_n725_c;
    logic fa_s0_c100_n726_s, fa_s0_c100_n726_c;
    logic fa_s0_c100_n727_s, fa_s0_c100_n727_c;
    logic fa_s0_c100_n728_s, fa_s0_c100_n728_c;
    logic fa_s0_c100_n729_s, fa_s0_c100_n729_c;
    logic fa_s0_c101_n730_s, fa_s0_c101_n730_c;
    logic fa_s0_c101_n731_s, fa_s0_c101_n731_c;
    logic fa_s0_c101_n732_s, fa_s0_c101_n732_c;
    logic fa_s0_c101_n733_s, fa_s0_c101_n733_c;
    logic fa_s0_c101_n734_s, fa_s0_c101_n734_c;
    logic fa_s0_c101_n735_s, fa_s0_c101_n735_c;
    logic fa_s0_c101_n736_s, fa_s0_c101_n736_c;
    logic fa_s0_c101_n737_s, fa_s0_c101_n737_c;
    logic fa_s0_c101_n738_s, fa_s0_c101_n738_c;
    logic fa_s0_c101_n739_s, fa_s0_c101_n739_c;
    logic fa_s0_c102_n740_s, fa_s0_c102_n740_c;
    logic fa_s0_c102_n741_s, fa_s0_c102_n741_c;
    logic fa_s0_c102_n742_s, fa_s0_c102_n742_c;
    logic fa_s0_c102_n743_s, fa_s0_c102_n743_c;
    logic fa_s0_c102_n744_s, fa_s0_c102_n744_c;
    logic fa_s0_c102_n745_s, fa_s0_c102_n745_c;
    logic fa_s0_c102_n746_s, fa_s0_c102_n746_c;
    logic fa_s0_c102_n747_s, fa_s0_c102_n747_c;
    logic fa_s0_c102_n748_s, fa_s0_c102_n748_c;
    logic fa_s0_c102_n749_s, fa_s0_c102_n749_c;
    logic fa_s0_c102_n750_s, fa_s0_c102_n750_c;
    logic fa_s0_c103_n751_s, fa_s0_c103_n751_c;
    logic fa_s0_c103_n752_s, fa_s0_c103_n752_c;
    logic fa_s0_c103_n753_s, fa_s0_c103_n753_c;
    logic fa_s0_c103_n754_s, fa_s0_c103_n754_c;
    logic fa_s0_c103_n755_s, fa_s0_c103_n755_c;
    logic fa_s0_c103_n756_s, fa_s0_c103_n756_c;
    logic fa_s0_c103_n757_s, fa_s0_c103_n757_c;
    logic fa_s0_c103_n758_s, fa_s0_c103_n758_c;
    logic fa_s0_c103_n759_s, fa_s0_c103_n759_c;
    logic fa_s0_c103_n760_s, fa_s0_c103_n760_c;
    logic fa_s0_c104_n761_s, fa_s0_c104_n761_c;
    logic fa_s0_c104_n762_s, fa_s0_c104_n762_c;
    logic fa_s0_c104_n763_s, fa_s0_c104_n763_c;
    logic fa_s0_c104_n764_s, fa_s0_c104_n764_c;
    logic fa_s0_c104_n765_s, fa_s0_c104_n765_c;
    logic fa_s0_c104_n766_s, fa_s0_c104_n766_c;
    logic fa_s0_c104_n767_s, fa_s0_c104_n767_c;
    logic fa_s0_c104_n768_s, fa_s0_c104_n768_c;
    logic fa_s0_c104_n769_s, fa_s0_c104_n769_c;
    logic fa_s0_c104_n770_s, fa_s0_c104_n770_c;
    logic fa_s0_c104_n771_s, fa_s0_c104_n771_c;
    logic fa_s0_c105_n772_s, fa_s0_c105_n772_c;
    logic fa_s0_c105_n773_s, fa_s0_c105_n773_c;
    logic fa_s0_c105_n774_s, fa_s0_c105_n774_c;
    logic fa_s0_c105_n775_s, fa_s0_c105_n775_c;
    logic fa_s0_c105_n776_s, fa_s0_c105_n776_c;
    logic fa_s0_c105_n777_s, fa_s0_c105_n777_c;
    logic fa_s0_c105_n778_s, fa_s0_c105_n778_c;
    logic fa_s0_c105_n779_s, fa_s0_c105_n779_c;
    logic fa_s0_c105_n780_s, fa_s0_c105_n780_c;
    logic fa_s0_c105_n781_s, fa_s0_c105_n781_c;
    logic fa_s0_c106_n782_s, fa_s0_c106_n782_c;
    logic fa_s0_c106_n783_s, fa_s0_c106_n783_c;
    logic fa_s0_c106_n784_s, fa_s0_c106_n784_c;
    logic fa_s0_c106_n785_s, fa_s0_c106_n785_c;
    logic fa_s0_c106_n786_s, fa_s0_c106_n786_c;
    logic fa_s0_c106_n787_s, fa_s0_c106_n787_c;
    logic fa_s0_c106_n788_s, fa_s0_c106_n788_c;
    logic fa_s0_c106_n789_s, fa_s0_c106_n789_c;
    logic fa_s0_c106_n790_s, fa_s0_c106_n790_c;
    logic fa_s0_c106_n791_s, fa_s0_c106_n791_c;
    logic fa_s0_c106_n792_s, fa_s0_c106_n792_c;
    logic fa_s0_c107_n793_s, fa_s0_c107_n793_c;
    logic fa_s0_c107_n794_s, fa_s0_c107_n794_c;
    logic fa_s0_c107_n795_s, fa_s0_c107_n795_c;
    logic fa_s0_c107_n796_s, fa_s0_c107_n796_c;
    logic fa_s0_c107_n797_s, fa_s0_c107_n797_c;
    logic fa_s0_c107_n798_s, fa_s0_c107_n798_c;
    logic fa_s0_c107_n799_s, fa_s0_c107_n799_c;
    logic fa_s0_c107_n800_s, fa_s0_c107_n800_c;
    logic fa_s0_c107_n801_s, fa_s0_c107_n801_c;
    logic fa_s0_c107_n802_s, fa_s0_c107_n802_c;
    logic fa_s0_c108_n803_s, fa_s0_c108_n803_c;
    logic fa_s0_c108_n804_s, fa_s0_c108_n804_c;
    logic fa_s0_c108_n805_s, fa_s0_c108_n805_c;
    logic fa_s0_c108_n806_s, fa_s0_c108_n806_c;
    logic fa_s0_c108_n807_s, fa_s0_c108_n807_c;
    logic fa_s0_c108_n808_s, fa_s0_c108_n808_c;
    logic fa_s0_c108_n809_s, fa_s0_c108_n809_c;
    logic fa_s0_c108_n810_s, fa_s0_c108_n810_c;
    logic fa_s0_c108_n811_s, fa_s0_c108_n811_c;
    logic fa_s0_c108_n812_s, fa_s0_c108_n812_c;
    logic fa_s0_c108_n813_s, fa_s0_c108_n813_c;
    logic fa_s0_c109_n814_s, fa_s0_c109_n814_c;
    logic fa_s0_c109_n815_s, fa_s0_c109_n815_c;
    logic fa_s0_c109_n816_s, fa_s0_c109_n816_c;
    logic fa_s0_c109_n817_s, fa_s0_c109_n817_c;
    logic fa_s0_c109_n818_s, fa_s0_c109_n818_c;
    logic fa_s0_c109_n819_s, fa_s0_c109_n819_c;
    logic fa_s0_c109_n820_s, fa_s0_c109_n820_c;
    logic fa_s0_c109_n821_s, fa_s0_c109_n821_c;
    logic fa_s0_c109_n822_s, fa_s0_c109_n822_c;
    logic fa_s0_c109_n823_s, fa_s0_c109_n823_c;
    logic fa_s0_c110_n824_s, fa_s0_c110_n824_c;
    logic fa_s0_c110_n825_s, fa_s0_c110_n825_c;
    logic fa_s0_c110_n826_s, fa_s0_c110_n826_c;
    logic fa_s0_c110_n827_s, fa_s0_c110_n827_c;
    logic fa_s0_c110_n828_s, fa_s0_c110_n828_c;
    logic fa_s0_c110_n829_s, fa_s0_c110_n829_c;
    logic fa_s0_c110_n830_s, fa_s0_c110_n830_c;
    logic fa_s0_c110_n831_s, fa_s0_c110_n831_c;
    logic fa_s0_c110_n832_s, fa_s0_c110_n832_c;
    logic fa_s0_c110_n833_s, fa_s0_c110_n833_c;
    logic fa_s0_c110_n834_s, fa_s0_c110_n834_c;
    logic fa_s0_c111_n835_s, fa_s0_c111_n835_c;
    logic fa_s0_c111_n836_s, fa_s0_c111_n836_c;
    logic fa_s0_c111_n837_s, fa_s0_c111_n837_c;
    logic fa_s0_c111_n838_s, fa_s0_c111_n838_c;
    logic fa_s0_c111_n839_s, fa_s0_c111_n839_c;
    logic fa_s0_c111_n840_s, fa_s0_c111_n840_c;
    logic fa_s0_c111_n841_s, fa_s0_c111_n841_c;
    logic fa_s0_c111_n842_s, fa_s0_c111_n842_c;
    logic fa_s0_c111_n843_s, fa_s0_c111_n843_c;
    logic fa_s0_c111_n844_s, fa_s0_c111_n844_c;
    logic fa_s0_c112_n845_s, fa_s0_c112_n845_c;
    logic fa_s0_c112_n846_s, fa_s0_c112_n846_c;
    logic fa_s0_c112_n847_s, fa_s0_c112_n847_c;
    logic fa_s0_c112_n848_s, fa_s0_c112_n848_c;
    logic fa_s0_c112_n849_s, fa_s0_c112_n849_c;
    logic fa_s0_c112_n850_s, fa_s0_c112_n850_c;
    logic fa_s0_c112_n851_s, fa_s0_c112_n851_c;
    logic fa_s0_c112_n852_s, fa_s0_c112_n852_c;
    logic fa_s0_c112_n853_s, fa_s0_c112_n853_c;
    logic fa_s0_c112_n854_s, fa_s0_c112_n854_c;
    logic fa_s0_c112_n855_s, fa_s0_c112_n855_c;
    logic fa_s0_c113_n856_s, fa_s0_c113_n856_c;
    logic fa_s0_c113_n857_s, fa_s0_c113_n857_c;
    logic fa_s0_c113_n858_s, fa_s0_c113_n858_c;
    logic fa_s0_c113_n859_s, fa_s0_c113_n859_c;
    logic fa_s0_c113_n860_s, fa_s0_c113_n860_c;
    logic fa_s0_c113_n861_s, fa_s0_c113_n861_c;
    logic fa_s0_c113_n862_s, fa_s0_c113_n862_c;
    logic fa_s0_c113_n863_s, fa_s0_c113_n863_c;
    logic fa_s0_c113_n864_s, fa_s0_c113_n864_c;
    logic fa_s0_c113_n865_s, fa_s0_c113_n865_c;
    logic fa_s0_c114_n866_s, fa_s0_c114_n866_c;
    logic fa_s0_c114_n867_s, fa_s0_c114_n867_c;
    logic fa_s0_c114_n868_s, fa_s0_c114_n868_c;
    logic fa_s0_c114_n869_s, fa_s0_c114_n869_c;
    logic fa_s0_c114_n870_s, fa_s0_c114_n870_c;
    logic fa_s0_c114_n871_s, fa_s0_c114_n871_c;
    logic fa_s0_c114_n872_s, fa_s0_c114_n872_c;
    logic fa_s0_c114_n873_s, fa_s0_c114_n873_c;
    logic fa_s0_c114_n874_s, fa_s0_c114_n874_c;
    logic fa_s0_c114_n875_s, fa_s0_c114_n875_c;
    logic fa_s0_c114_n876_s, fa_s0_c114_n876_c;
    logic fa_s0_c115_n877_s, fa_s0_c115_n877_c;
    logic fa_s0_c115_n878_s, fa_s0_c115_n878_c;
    logic fa_s0_c115_n879_s, fa_s0_c115_n879_c;
    logic fa_s0_c115_n880_s, fa_s0_c115_n880_c;
    logic fa_s0_c115_n881_s, fa_s0_c115_n881_c;
    logic fa_s0_c115_n882_s, fa_s0_c115_n882_c;
    logic fa_s0_c115_n883_s, fa_s0_c115_n883_c;
    logic fa_s0_c115_n884_s, fa_s0_c115_n884_c;
    logic fa_s0_c115_n885_s, fa_s0_c115_n885_c;
    logic fa_s0_c115_n886_s, fa_s0_c115_n886_c;
    logic fa_s0_c116_n887_s, fa_s0_c116_n887_c;
    logic fa_s0_c116_n888_s, fa_s0_c116_n888_c;
    logic fa_s0_c116_n889_s, fa_s0_c116_n889_c;
    logic fa_s0_c116_n890_s, fa_s0_c116_n890_c;
    logic fa_s0_c116_n891_s, fa_s0_c116_n891_c;
    logic fa_s0_c116_n892_s, fa_s0_c116_n892_c;
    logic fa_s0_c116_n893_s, fa_s0_c116_n893_c;
    logic fa_s0_c116_n894_s, fa_s0_c116_n894_c;
    logic fa_s0_c116_n895_s, fa_s0_c116_n895_c;
    logic fa_s0_c116_n896_s, fa_s0_c116_n896_c;
    logic fa_s0_c116_n897_s, fa_s0_c116_n897_c;
    logic fa_s0_c117_n898_s, fa_s0_c117_n898_c;
    logic fa_s0_c117_n899_s, fa_s0_c117_n899_c;
    logic fa_s0_c117_n900_s, fa_s0_c117_n900_c;
    logic fa_s0_c117_n901_s, fa_s0_c117_n901_c;
    logic fa_s0_c117_n902_s, fa_s0_c117_n902_c;
    logic fa_s0_c117_n903_s, fa_s0_c117_n903_c;
    logic fa_s0_c117_n904_s, fa_s0_c117_n904_c;
    logic fa_s0_c117_n905_s, fa_s0_c117_n905_c;
    logic fa_s0_c117_n906_s, fa_s0_c117_n906_c;
    logic fa_s0_c117_n907_s, fa_s0_c117_n907_c;
    logic fa_s0_c118_n908_s, fa_s0_c118_n908_c;
    logic fa_s0_c118_n909_s, fa_s0_c118_n909_c;
    logic fa_s0_c118_n910_s, fa_s0_c118_n910_c;
    logic fa_s0_c118_n911_s, fa_s0_c118_n911_c;
    logic fa_s0_c118_n912_s, fa_s0_c118_n912_c;
    logic fa_s0_c118_n913_s, fa_s0_c118_n913_c;
    logic fa_s0_c118_n914_s, fa_s0_c118_n914_c;
    logic fa_s0_c118_n915_s, fa_s0_c118_n915_c;
    logic fa_s0_c118_n916_s, fa_s0_c118_n916_c;
    logic fa_s0_c118_n917_s, fa_s0_c118_n917_c;
    logic fa_s0_c118_n918_s, fa_s0_c118_n918_c;
    logic fa_s0_c119_n919_s, fa_s0_c119_n919_c;
    logic fa_s0_c119_n920_s, fa_s0_c119_n920_c;
    logic fa_s0_c119_n921_s, fa_s0_c119_n921_c;
    logic fa_s0_c119_n922_s, fa_s0_c119_n922_c;
    logic fa_s0_c119_n923_s, fa_s0_c119_n923_c;
    logic fa_s0_c119_n924_s, fa_s0_c119_n924_c;
    logic fa_s0_c119_n925_s, fa_s0_c119_n925_c;
    logic fa_s0_c119_n926_s, fa_s0_c119_n926_c;
    logic fa_s0_c119_n927_s, fa_s0_c119_n927_c;
    logic fa_s0_c119_n928_s, fa_s0_c119_n928_c;
    logic fa_s0_c120_n929_s, fa_s0_c120_n929_c;
    logic fa_s0_c120_n930_s, fa_s0_c120_n930_c;
    logic fa_s0_c120_n931_s, fa_s0_c120_n931_c;
    logic fa_s0_c120_n932_s, fa_s0_c120_n932_c;
    logic fa_s0_c120_n933_s, fa_s0_c120_n933_c;
    logic fa_s0_c120_n934_s, fa_s0_c120_n934_c;
    logic fa_s0_c120_n935_s, fa_s0_c120_n935_c;
    logic fa_s0_c120_n936_s, fa_s0_c120_n936_c;
    logic fa_s0_c120_n937_s, fa_s0_c120_n937_c;
    logic fa_s0_c120_n938_s, fa_s0_c120_n938_c;
    logic fa_s0_c120_n939_s, fa_s0_c120_n939_c;
    logic fa_s0_c121_n940_s, fa_s0_c121_n940_c;
    logic fa_s0_c121_n941_s, fa_s0_c121_n941_c;
    logic fa_s0_c121_n942_s, fa_s0_c121_n942_c;
    logic fa_s0_c121_n943_s, fa_s0_c121_n943_c;
    logic fa_s0_c121_n944_s, fa_s0_c121_n944_c;
    logic fa_s0_c121_n945_s, fa_s0_c121_n945_c;
    logic fa_s0_c121_n946_s, fa_s0_c121_n946_c;
    logic fa_s0_c121_n947_s, fa_s0_c121_n947_c;
    logic fa_s0_c121_n948_s, fa_s0_c121_n948_c;
    logic fa_s0_c121_n949_s, fa_s0_c121_n949_c;
    logic fa_s0_c122_n950_s, fa_s0_c122_n950_c;
    logic fa_s0_c122_n951_s, fa_s0_c122_n951_c;
    logic fa_s0_c122_n952_s, fa_s0_c122_n952_c;
    logic fa_s0_c122_n953_s, fa_s0_c122_n953_c;
    logic fa_s0_c122_n954_s, fa_s0_c122_n954_c;
    logic fa_s0_c122_n955_s, fa_s0_c122_n955_c;
    logic fa_s0_c122_n956_s, fa_s0_c122_n956_c;
    logic fa_s0_c122_n957_s, fa_s0_c122_n957_c;
    logic fa_s0_c122_n958_s, fa_s0_c122_n958_c;
    logic fa_s0_c122_n959_s, fa_s0_c122_n959_c;
    logic fa_s0_c122_n960_s, fa_s0_c122_n960_c;
    logic fa_s0_c123_n961_s, fa_s0_c123_n961_c;
    logic fa_s0_c123_n962_s, fa_s0_c123_n962_c;
    logic fa_s0_c123_n963_s, fa_s0_c123_n963_c;
    logic fa_s0_c123_n964_s, fa_s0_c123_n964_c;
    logic fa_s0_c123_n965_s, fa_s0_c123_n965_c;
    logic fa_s0_c123_n966_s, fa_s0_c123_n966_c;
    logic fa_s0_c123_n967_s, fa_s0_c123_n967_c;
    logic fa_s0_c123_n968_s, fa_s0_c123_n968_c;
    logic fa_s0_c123_n969_s, fa_s0_c123_n969_c;
    logic fa_s0_c123_n970_s, fa_s0_c123_n970_c;
    logic fa_s0_c124_n971_s, fa_s0_c124_n971_c;
    logic fa_s0_c124_n972_s, fa_s0_c124_n972_c;
    logic fa_s0_c124_n973_s, fa_s0_c124_n973_c;
    logic fa_s0_c124_n974_s, fa_s0_c124_n974_c;
    logic fa_s0_c124_n975_s, fa_s0_c124_n975_c;
    logic fa_s0_c124_n976_s, fa_s0_c124_n976_c;
    logic fa_s0_c124_n977_s, fa_s0_c124_n977_c;
    logic fa_s0_c124_n978_s, fa_s0_c124_n978_c;
    logic fa_s0_c124_n979_s, fa_s0_c124_n979_c;
    logic fa_s0_c124_n980_s, fa_s0_c124_n980_c;
    logic fa_s0_c124_n981_s, fa_s0_c124_n981_c;
    logic fa_s0_c125_n982_s, fa_s0_c125_n982_c;
    logic fa_s0_c125_n983_s, fa_s0_c125_n983_c;
    logic fa_s0_c125_n984_s, fa_s0_c125_n984_c;
    logic fa_s0_c125_n985_s, fa_s0_c125_n985_c;
    logic fa_s0_c125_n986_s, fa_s0_c125_n986_c;
    logic fa_s0_c125_n987_s, fa_s0_c125_n987_c;
    logic fa_s0_c125_n988_s, fa_s0_c125_n988_c;
    logic fa_s0_c125_n989_s, fa_s0_c125_n989_c;
    logic fa_s0_c125_n990_s, fa_s0_c125_n990_c;
    logic fa_s0_c125_n991_s, fa_s0_c125_n991_c;
    logic fa_s0_c126_n992_s, fa_s0_c126_n992_c;
    logic fa_s0_c126_n993_s, fa_s0_c126_n993_c;
    logic fa_s0_c126_n994_s, fa_s0_c126_n994_c;
    logic fa_s0_c126_n995_s, fa_s0_c126_n995_c;
    logic fa_s0_c126_n996_s, fa_s0_c126_n996_c;
    logic fa_s0_c126_n997_s, fa_s0_c126_n997_c;
    logic fa_s0_c126_n998_s, fa_s0_c126_n998_c;
    logic fa_s0_c126_n999_s, fa_s0_c126_n999_c;
    logic fa_s0_c126_n1000_s, fa_s0_c126_n1000_c;
    logic fa_s0_c126_n1001_s, fa_s0_c126_n1001_c;
    logic fa_s0_c126_n1002_s, fa_s0_c126_n1002_c;
    logic fa_s1_c3_n0_s, fa_s1_c3_n0_c;
    logic fa_s1_c6_n1_s, fa_s1_c6_n1_c;
    logic fa_s1_c7_n2_s, fa_s1_c7_n2_c;
    logic fa_s1_c8_n3_s, fa_s1_c8_n3_c;
    logic fa_s1_c9_n4_s, fa_s1_c9_n4_c;
    logic fa_s1_c10_n5_s, fa_s1_c10_n5_c;
    logic fa_s1_c11_n6_s, fa_s1_c11_n6_c;
    logic fa_s1_c12_n7_s, fa_s1_c12_n7_c;
    logic fa_s1_c12_n8_s, fa_s1_c12_n8_c;
    logic fa_s1_c13_n9_s, fa_s1_c13_n9_c;
    logic fa_s1_c14_n10_s, fa_s1_c14_n10_c;
    logic fa_s1_c15_n11_s, fa_s1_c15_n11_c;
    logic fa_s1_c15_n12_s, fa_s1_c15_n12_c;
    logic fa_s1_c16_n13_s, fa_s1_c16_n13_c;
    logic fa_s1_c16_n14_s, fa_s1_c16_n14_c;
    logic fa_s1_c17_n15_s, fa_s1_c17_n15_c;
    logic fa_s1_c17_n16_s, fa_s1_c17_n16_c;
    logic fa_s1_c18_n17_s, fa_s1_c18_n17_c;
    logic fa_s1_c18_n18_s, fa_s1_c18_n18_c;
    logic fa_s1_c19_n19_s, fa_s1_c19_n19_c;
    logic fa_s1_c19_n20_s, fa_s1_c19_n20_c;
    logic fa_s1_c20_n21_s, fa_s1_c20_n21_c;
    logic fa_s1_c20_n22_s, fa_s1_c20_n22_c;
    logic fa_s1_c21_n23_s, fa_s1_c21_n23_c;
    logic fa_s1_c21_n24_s, fa_s1_c21_n24_c;
    logic fa_s1_c21_n25_s, fa_s1_c21_n25_c;
    logic fa_s1_c22_n26_s, fa_s1_c22_n26_c;
    logic fa_s1_c22_n27_s, fa_s1_c22_n27_c;
    logic fa_s1_c23_n28_s, fa_s1_c23_n28_c;
    logic fa_s1_c23_n29_s, fa_s1_c23_n29_c;
    logic fa_s1_c24_n30_s, fa_s1_c24_n30_c;
    logic fa_s1_c24_n31_s, fa_s1_c24_n31_c;
    logic fa_s1_c24_n32_s, fa_s1_c24_n32_c;
    logic fa_s1_c25_n33_s, fa_s1_c25_n33_c;
    logic fa_s1_c25_n34_s, fa_s1_c25_n34_c;
    logic fa_s1_c25_n35_s, fa_s1_c25_n35_c;
    logic fa_s1_c26_n36_s, fa_s1_c26_n36_c;
    logic fa_s1_c26_n37_s, fa_s1_c26_n37_c;
    logic fa_s1_c26_n38_s, fa_s1_c26_n38_c;
    logic fa_s1_c27_n39_s, fa_s1_c27_n39_c;
    logic fa_s1_c27_n40_s, fa_s1_c27_n40_c;
    logic fa_s1_c27_n41_s, fa_s1_c27_n41_c;
    logic fa_s1_c28_n42_s, fa_s1_c28_n42_c;
    logic fa_s1_c28_n43_s, fa_s1_c28_n43_c;
    logic fa_s1_c28_n44_s, fa_s1_c28_n44_c;
    logic fa_s1_c29_n45_s, fa_s1_c29_n45_c;
    logic fa_s1_c29_n46_s, fa_s1_c29_n46_c;
    logic fa_s1_c29_n47_s, fa_s1_c29_n47_c;
    logic fa_s1_c30_n48_s, fa_s1_c30_n48_c;
    logic fa_s1_c30_n49_s, fa_s1_c30_n49_c;
    logic fa_s1_c30_n50_s, fa_s1_c30_n50_c;
    logic fa_s1_c30_n51_s, fa_s1_c30_n51_c;
    logic fa_s1_c31_n52_s, fa_s1_c31_n52_c;
    logic fa_s1_c31_n53_s, fa_s1_c31_n53_c;
    logic fa_s1_c31_n54_s, fa_s1_c31_n54_c;
    logic fa_s1_c32_n55_s, fa_s1_c32_n55_c;
    logic fa_s1_c32_n56_s, fa_s1_c32_n56_c;
    logic fa_s1_c32_n57_s, fa_s1_c32_n57_c;
    logic fa_s1_c33_n58_s, fa_s1_c33_n58_c;
    logic fa_s1_c33_n59_s, fa_s1_c33_n59_c;
    logic fa_s1_c33_n60_s, fa_s1_c33_n60_c;
    logic fa_s1_c33_n61_s, fa_s1_c33_n61_c;
    logic fa_s1_c34_n62_s, fa_s1_c34_n62_c;
    logic fa_s1_c34_n63_s, fa_s1_c34_n63_c;
    logic fa_s1_c34_n64_s, fa_s1_c34_n64_c;
    logic fa_s1_c34_n65_s, fa_s1_c34_n65_c;
    logic fa_s1_c35_n66_s, fa_s1_c35_n66_c;
    logic fa_s1_c35_n67_s, fa_s1_c35_n67_c;
    logic fa_s1_c35_n68_s, fa_s1_c35_n68_c;
    logic fa_s1_c35_n69_s, fa_s1_c35_n69_c;
    logic fa_s1_c36_n70_s, fa_s1_c36_n70_c;
    logic fa_s1_c36_n71_s, fa_s1_c36_n71_c;
    logic fa_s1_c36_n72_s, fa_s1_c36_n72_c;
    logic fa_s1_c36_n73_s, fa_s1_c36_n73_c;
    logic fa_s1_c37_n74_s, fa_s1_c37_n74_c;
    logic fa_s1_c37_n75_s, fa_s1_c37_n75_c;
    logic fa_s1_c37_n76_s, fa_s1_c37_n76_c;
    logic fa_s1_c37_n77_s, fa_s1_c37_n77_c;
    logic fa_s1_c38_n78_s, fa_s1_c38_n78_c;
    logic fa_s1_c38_n79_s, fa_s1_c38_n79_c;
    logic fa_s1_c38_n80_s, fa_s1_c38_n80_c;
    logic fa_s1_c38_n81_s, fa_s1_c38_n81_c;
    logic fa_s1_c39_n82_s, fa_s1_c39_n82_c;
    logic fa_s1_c39_n83_s, fa_s1_c39_n83_c;
    logic fa_s1_c39_n84_s, fa_s1_c39_n84_c;
    logic fa_s1_c39_n85_s, fa_s1_c39_n85_c;
    logic fa_s1_c39_n86_s, fa_s1_c39_n86_c;
    logic fa_s1_c40_n87_s, fa_s1_c40_n87_c;
    logic fa_s1_c40_n88_s, fa_s1_c40_n88_c;
    logic fa_s1_c40_n89_s, fa_s1_c40_n89_c;
    logic fa_s1_c40_n90_s, fa_s1_c40_n90_c;
    logic fa_s1_c41_n91_s, fa_s1_c41_n91_c;
    logic fa_s1_c41_n92_s, fa_s1_c41_n92_c;
    logic fa_s1_c41_n93_s, fa_s1_c41_n93_c;
    logic fa_s1_c41_n94_s, fa_s1_c41_n94_c;
    logic fa_s1_c42_n95_s, fa_s1_c42_n95_c;
    logic fa_s1_c42_n96_s, fa_s1_c42_n96_c;
    logic fa_s1_c42_n97_s, fa_s1_c42_n97_c;
    logic fa_s1_c42_n98_s, fa_s1_c42_n98_c;
    logic fa_s1_c42_n99_s, fa_s1_c42_n99_c;
    logic fa_s1_c43_n100_s, fa_s1_c43_n100_c;
    logic fa_s1_c43_n101_s, fa_s1_c43_n101_c;
    logic fa_s1_c43_n102_s, fa_s1_c43_n102_c;
    logic fa_s1_c43_n103_s, fa_s1_c43_n103_c;
    logic fa_s1_c43_n104_s, fa_s1_c43_n104_c;
    logic fa_s1_c44_n105_s, fa_s1_c44_n105_c;
    logic fa_s1_c44_n106_s, fa_s1_c44_n106_c;
    logic fa_s1_c44_n107_s, fa_s1_c44_n107_c;
    logic fa_s1_c44_n108_s, fa_s1_c44_n108_c;
    logic fa_s1_c44_n109_s, fa_s1_c44_n109_c;
    logic fa_s1_c45_n110_s, fa_s1_c45_n110_c;
    logic fa_s1_c45_n111_s, fa_s1_c45_n111_c;
    logic fa_s1_c45_n112_s, fa_s1_c45_n112_c;
    logic fa_s1_c45_n113_s, fa_s1_c45_n113_c;
    logic fa_s1_c45_n114_s, fa_s1_c45_n114_c;
    logic fa_s1_c46_n115_s, fa_s1_c46_n115_c;
    logic fa_s1_c46_n116_s, fa_s1_c46_n116_c;
    logic fa_s1_c46_n117_s, fa_s1_c46_n117_c;
    logic fa_s1_c46_n118_s, fa_s1_c46_n118_c;
    logic fa_s1_c46_n119_s, fa_s1_c46_n119_c;
    logic fa_s1_c47_n120_s, fa_s1_c47_n120_c;
    logic fa_s1_c47_n121_s, fa_s1_c47_n121_c;
    logic fa_s1_c47_n122_s, fa_s1_c47_n122_c;
    logic fa_s1_c47_n123_s, fa_s1_c47_n123_c;
    logic fa_s1_c47_n124_s, fa_s1_c47_n124_c;
    logic fa_s1_c48_n125_s, fa_s1_c48_n125_c;
    logic fa_s1_c48_n126_s, fa_s1_c48_n126_c;
    logic fa_s1_c48_n127_s, fa_s1_c48_n127_c;
    logic fa_s1_c48_n128_s, fa_s1_c48_n128_c;
    logic fa_s1_c48_n129_s, fa_s1_c48_n129_c;
    logic fa_s1_c48_n130_s, fa_s1_c48_n130_c;
    logic fa_s1_c49_n131_s, fa_s1_c49_n131_c;
    logic fa_s1_c49_n132_s, fa_s1_c49_n132_c;
    logic fa_s1_c49_n133_s, fa_s1_c49_n133_c;
    logic fa_s1_c49_n134_s, fa_s1_c49_n134_c;
    logic fa_s1_c49_n135_s, fa_s1_c49_n135_c;
    logic fa_s1_c50_n136_s, fa_s1_c50_n136_c;
    logic fa_s1_c50_n137_s, fa_s1_c50_n137_c;
    logic fa_s1_c50_n138_s, fa_s1_c50_n138_c;
    logic fa_s1_c50_n139_s, fa_s1_c50_n139_c;
    logic fa_s1_c50_n140_s, fa_s1_c50_n140_c;
    logic fa_s1_c51_n141_s, fa_s1_c51_n141_c;
    logic fa_s1_c51_n142_s, fa_s1_c51_n142_c;
    logic fa_s1_c51_n143_s, fa_s1_c51_n143_c;
    logic fa_s1_c51_n144_s, fa_s1_c51_n144_c;
    logic fa_s1_c51_n145_s, fa_s1_c51_n145_c;
    logic fa_s1_c51_n146_s, fa_s1_c51_n146_c;
    logic fa_s1_c52_n147_s, fa_s1_c52_n147_c;
    logic fa_s1_c52_n148_s, fa_s1_c52_n148_c;
    logic fa_s1_c52_n149_s, fa_s1_c52_n149_c;
    logic fa_s1_c52_n150_s, fa_s1_c52_n150_c;
    logic fa_s1_c52_n151_s, fa_s1_c52_n151_c;
    logic fa_s1_c52_n152_s, fa_s1_c52_n152_c;
    logic fa_s1_c53_n153_s, fa_s1_c53_n153_c;
    logic fa_s1_c53_n154_s, fa_s1_c53_n154_c;
    logic fa_s1_c53_n155_s, fa_s1_c53_n155_c;
    logic fa_s1_c53_n156_s, fa_s1_c53_n156_c;
    logic fa_s1_c53_n157_s, fa_s1_c53_n157_c;
    logic fa_s1_c53_n158_s, fa_s1_c53_n158_c;
    logic fa_s1_c54_n159_s, fa_s1_c54_n159_c;
    logic fa_s1_c54_n160_s, fa_s1_c54_n160_c;
    logic fa_s1_c54_n161_s, fa_s1_c54_n161_c;
    logic fa_s1_c54_n162_s, fa_s1_c54_n162_c;
    logic fa_s1_c54_n163_s, fa_s1_c54_n163_c;
    logic fa_s1_c54_n164_s, fa_s1_c54_n164_c;
    logic fa_s1_c55_n165_s, fa_s1_c55_n165_c;
    logic fa_s1_c55_n166_s, fa_s1_c55_n166_c;
    logic fa_s1_c55_n167_s, fa_s1_c55_n167_c;
    logic fa_s1_c55_n168_s, fa_s1_c55_n168_c;
    logic fa_s1_c55_n169_s, fa_s1_c55_n169_c;
    logic fa_s1_c55_n170_s, fa_s1_c55_n170_c;
    logic fa_s1_c56_n171_s, fa_s1_c56_n171_c;
    logic fa_s1_c56_n172_s, fa_s1_c56_n172_c;
    logic fa_s1_c56_n173_s, fa_s1_c56_n173_c;
    logic fa_s1_c56_n174_s, fa_s1_c56_n174_c;
    logic fa_s1_c56_n175_s, fa_s1_c56_n175_c;
    logic fa_s1_c56_n176_s, fa_s1_c56_n176_c;
    logic fa_s1_c57_n177_s, fa_s1_c57_n177_c;
    logic fa_s1_c57_n178_s, fa_s1_c57_n178_c;
    logic fa_s1_c57_n179_s, fa_s1_c57_n179_c;
    logic fa_s1_c57_n180_s, fa_s1_c57_n180_c;
    logic fa_s1_c57_n181_s, fa_s1_c57_n181_c;
    logic fa_s1_c57_n182_s, fa_s1_c57_n182_c;
    logic fa_s1_c57_n183_s, fa_s1_c57_n183_c;
    logic fa_s1_c58_n184_s, fa_s1_c58_n184_c;
    logic fa_s1_c58_n185_s, fa_s1_c58_n185_c;
    logic fa_s1_c58_n186_s, fa_s1_c58_n186_c;
    logic fa_s1_c58_n187_s, fa_s1_c58_n187_c;
    logic fa_s1_c58_n188_s, fa_s1_c58_n188_c;
    logic fa_s1_c58_n189_s, fa_s1_c58_n189_c;
    logic fa_s1_c59_n190_s, fa_s1_c59_n190_c;
    logic fa_s1_c59_n191_s, fa_s1_c59_n191_c;
    logic fa_s1_c59_n192_s, fa_s1_c59_n192_c;
    logic fa_s1_c59_n193_s, fa_s1_c59_n193_c;
    logic fa_s1_c59_n194_s, fa_s1_c59_n194_c;
    logic fa_s1_c59_n195_s, fa_s1_c59_n195_c;
    logic fa_s1_c60_n196_s, fa_s1_c60_n196_c;
    logic fa_s1_c60_n197_s, fa_s1_c60_n197_c;
    logic fa_s1_c60_n198_s, fa_s1_c60_n198_c;
    logic fa_s1_c60_n199_s, fa_s1_c60_n199_c;
    logic fa_s1_c60_n200_s, fa_s1_c60_n200_c;
    logic fa_s1_c60_n201_s, fa_s1_c60_n201_c;
    logic fa_s1_c60_n202_s, fa_s1_c60_n202_c;
    logic fa_s1_c61_n203_s, fa_s1_c61_n203_c;
    logic fa_s1_c61_n204_s, fa_s1_c61_n204_c;
    logic fa_s1_c61_n205_s, fa_s1_c61_n205_c;
    logic fa_s1_c61_n206_s, fa_s1_c61_n206_c;
    logic fa_s1_c61_n207_s, fa_s1_c61_n207_c;
    logic fa_s1_c61_n208_s, fa_s1_c61_n208_c;
    logic fa_s1_c61_n209_s, fa_s1_c61_n209_c;
    logic fa_s1_c62_n210_s, fa_s1_c62_n210_c;
    logic fa_s1_c62_n211_s, fa_s1_c62_n211_c;
    logic fa_s1_c62_n212_s, fa_s1_c62_n212_c;
    logic fa_s1_c62_n213_s, fa_s1_c62_n213_c;
    logic fa_s1_c62_n214_s, fa_s1_c62_n214_c;
    logic fa_s1_c62_n215_s, fa_s1_c62_n215_c;
    logic fa_s1_c62_n216_s, fa_s1_c62_n216_c;
    logic fa_s1_c63_n217_s, fa_s1_c63_n217_c;
    logic fa_s1_c63_n218_s, fa_s1_c63_n218_c;
    logic fa_s1_c63_n219_s, fa_s1_c63_n219_c;
    logic fa_s1_c63_n220_s, fa_s1_c63_n220_c;
    logic fa_s1_c63_n221_s, fa_s1_c63_n221_c;
    logic fa_s1_c63_n222_s, fa_s1_c63_n222_c;
    logic fa_s1_c63_n223_s, fa_s1_c63_n223_c;
    logic fa_s1_c64_n224_s, fa_s1_c64_n224_c;
    logic fa_s1_c64_n225_s, fa_s1_c64_n225_c;
    logic fa_s1_c64_n226_s, fa_s1_c64_n226_c;
    logic fa_s1_c64_n227_s, fa_s1_c64_n227_c;
    logic fa_s1_c64_n228_s, fa_s1_c64_n228_c;
    logic fa_s1_c64_n229_s, fa_s1_c64_n229_c;
    logic fa_s1_c64_n230_s, fa_s1_c64_n230_c;
    logic fa_s1_c65_n231_s, fa_s1_c65_n231_c;
    logic fa_s1_c65_n232_s, fa_s1_c65_n232_c;
    logic fa_s1_c65_n233_s, fa_s1_c65_n233_c;
    logic fa_s1_c65_n234_s, fa_s1_c65_n234_c;
    logic fa_s1_c65_n235_s, fa_s1_c65_n235_c;
    logic fa_s1_c65_n236_s, fa_s1_c65_n236_c;
    logic fa_s1_c65_n237_s, fa_s1_c65_n237_c;
    logic fa_s1_c66_n238_s, fa_s1_c66_n238_c;
    logic fa_s1_c66_n239_s, fa_s1_c66_n239_c;
    logic fa_s1_c66_n240_s, fa_s1_c66_n240_c;
    logic fa_s1_c66_n241_s, fa_s1_c66_n241_c;
    logic fa_s1_c66_n242_s, fa_s1_c66_n242_c;
    logic fa_s1_c66_n243_s, fa_s1_c66_n243_c;
    logic fa_s1_c66_n244_s, fa_s1_c66_n244_c;
    logic fa_s1_c67_n245_s, fa_s1_c67_n245_c;
    logic fa_s1_c67_n246_s, fa_s1_c67_n246_c;
    logic fa_s1_c67_n247_s, fa_s1_c67_n247_c;
    logic fa_s1_c67_n248_s, fa_s1_c67_n248_c;
    logic fa_s1_c67_n249_s, fa_s1_c67_n249_c;
    logic fa_s1_c67_n250_s, fa_s1_c67_n250_c;
    logic fa_s1_c67_n251_s, fa_s1_c67_n251_c;
    logic fa_s1_c68_n252_s, fa_s1_c68_n252_c;
    logic fa_s1_c68_n253_s, fa_s1_c68_n253_c;
    logic fa_s1_c68_n254_s, fa_s1_c68_n254_c;
    logic fa_s1_c68_n255_s, fa_s1_c68_n255_c;
    logic fa_s1_c68_n256_s, fa_s1_c68_n256_c;
    logic fa_s1_c68_n257_s, fa_s1_c68_n257_c;
    logic fa_s1_c68_n258_s, fa_s1_c68_n258_c;
    logic fa_s1_c69_n259_s, fa_s1_c69_n259_c;
    logic fa_s1_c69_n260_s, fa_s1_c69_n260_c;
    logic fa_s1_c69_n261_s, fa_s1_c69_n261_c;
    logic fa_s1_c69_n262_s, fa_s1_c69_n262_c;
    logic fa_s1_c69_n263_s, fa_s1_c69_n263_c;
    logic fa_s1_c69_n264_s, fa_s1_c69_n264_c;
    logic fa_s1_c69_n265_s, fa_s1_c69_n265_c;
    logic fa_s1_c70_n266_s, fa_s1_c70_n266_c;
    logic fa_s1_c70_n267_s, fa_s1_c70_n267_c;
    logic fa_s1_c70_n268_s, fa_s1_c70_n268_c;
    logic fa_s1_c70_n269_s, fa_s1_c70_n269_c;
    logic fa_s1_c70_n270_s, fa_s1_c70_n270_c;
    logic fa_s1_c70_n271_s, fa_s1_c70_n271_c;
    logic fa_s1_c70_n272_s, fa_s1_c70_n272_c;
    logic fa_s1_c71_n273_s, fa_s1_c71_n273_c;
    logic fa_s1_c71_n274_s, fa_s1_c71_n274_c;
    logic fa_s1_c71_n275_s, fa_s1_c71_n275_c;
    logic fa_s1_c71_n276_s, fa_s1_c71_n276_c;
    logic fa_s1_c71_n277_s, fa_s1_c71_n277_c;
    logic fa_s1_c71_n278_s, fa_s1_c71_n278_c;
    logic fa_s1_c71_n279_s, fa_s1_c71_n279_c;
    logic fa_s1_c72_n280_s, fa_s1_c72_n280_c;
    logic fa_s1_c72_n281_s, fa_s1_c72_n281_c;
    logic fa_s1_c72_n282_s, fa_s1_c72_n282_c;
    logic fa_s1_c72_n283_s, fa_s1_c72_n283_c;
    logic fa_s1_c72_n284_s, fa_s1_c72_n284_c;
    logic fa_s1_c72_n285_s, fa_s1_c72_n285_c;
    logic fa_s1_c72_n286_s, fa_s1_c72_n286_c;
    logic fa_s1_c73_n287_s, fa_s1_c73_n287_c;
    logic fa_s1_c73_n288_s, fa_s1_c73_n288_c;
    logic fa_s1_c73_n289_s, fa_s1_c73_n289_c;
    logic fa_s1_c73_n290_s, fa_s1_c73_n290_c;
    logic fa_s1_c73_n291_s, fa_s1_c73_n291_c;
    logic fa_s1_c73_n292_s, fa_s1_c73_n292_c;
    logic fa_s1_c73_n293_s, fa_s1_c73_n293_c;
    logic fa_s1_c74_n294_s, fa_s1_c74_n294_c;
    logic fa_s1_c74_n295_s, fa_s1_c74_n295_c;
    logic fa_s1_c74_n296_s, fa_s1_c74_n296_c;
    logic fa_s1_c74_n297_s, fa_s1_c74_n297_c;
    logic fa_s1_c74_n298_s, fa_s1_c74_n298_c;
    logic fa_s1_c74_n299_s, fa_s1_c74_n299_c;
    logic fa_s1_c74_n300_s, fa_s1_c74_n300_c;
    logic fa_s1_c75_n301_s, fa_s1_c75_n301_c;
    logic fa_s1_c75_n302_s, fa_s1_c75_n302_c;
    logic fa_s1_c75_n303_s, fa_s1_c75_n303_c;
    logic fa_s1_c75_n304_s, fa_s1_c75_n304_c;
    logic fa_s1_c75_n305_s, fa_s1_c75_n305_c;
    logic fa_s1_c75_n306_s, fa_s1_c75_n306_c;
    logic fa_s1_c75_n307_s, fa_s1_c75_n307_c;
    logic fa_s1_c76_n308_s, fa_s1_c76_n308_c;
    logic fa_s1_c76_n309_s, fa_s1_c76_n309_c;
    logic fa_s1_c76_n310_s, fa_s1_c76_n310_c;
    logic fa_s1_c76_n311_s, fa_s1_c76_n311_c;
    logic fa_s1_c76_n312_s, fa_s1_c76_n312_c;
    logic fa_s1_c76_n313_s, fa_s1_c76_n313_c;
    logic fa_s1_c76_n314_s, fa_s1_c76_n314_c;
    logic fa_s1_c77_n315_s, fa_s1_c77_n315_c;
    logic fa_s1_c77_n316_s, fa_s1_c77_n316_c;
    logic fa_s1_c77_n317_s, fa_s1_c77_n317_c;
    logic fa_s1_c77_n318_s, fa_s1_c77_n318_c;
    logic fa_s1_c77_n319_s, fa_s1_c77_n319_c;
    logic fa_s1_c77_n320_s, fa_s1_c77_n320_c;
    logic fa_s1_c77_n321_s, fa_s1_c77_n321_c;
    logic fa_s1_c78_n322_s, fa_s1_c78_n322_c;
    logic fa_s1_c78_n323_s, fa_s1_c78_n323_c;
    logic fa_s1_c78_n324_s, fa_s1_c78_n324_c;
    logic fa_s1_c78_n325_s, fa_s1_c78_n325_c;
    logic fa_s1_c78_n326_s, fa_s1_c78_n326_c;
    logic fa_s1_c78_n327_s, fa_s1_c78_n327_c;
    logic fa_s1_c78_n328_s, fa_s1_c78_n328_c;
    logic fa_s1_c79_n329_s, fa_s1_c79_n329_c;
    logic fa_s1_c79_n330_s, fa_s1_c79_n330_c;
    logic fa_s1_c79_n331_s, fa_s1_c79_n331_c;
    logic fa_s1_c79_n332_s, fa_s1_c79_n332_c;
    logic fa_s1_c79_n333_s, fa_s1_c79_n333_c;
    logic fa_s1_c79_n334_s, fa_s1_c79_n334_c;
    logic fa_s1_c79_n335_s, fa_s1_c79_n335_c;
    logic fa_s1_c80_n336_s, fa_s1_c80_n336_c;
    logic fa_s1_c80_n337_s, fa_s1_c80_n337_c;
    logic fa_s1_c80_n338_s, fa_s1_c80_n338_c;
    logic fa_s1_c80_n339_s, fa_s1_c80_n339_c;
    logic fa_s1_c80_n340_s, fa_s1_c80_n340_c;
    logic fa_s1_c80_n341_s, fa_s1_c80_n341_c;
    logic fa_s1_c80_n342_s, fa_s1_c80_n342_c;
    logic fa_s1_c81_n343_s, fa_s1_c81_n343_c;
    logic fa_s1_c81_n344_s, fa_s1_c81_n344_c;
    logic fa_s1_c81_n345_s, fa_s1_c81_n345_c;
    logic fa_s1_c81_n346_s, fa_s1_c81_n346_c;
    logic fa_s1_c81_n347_s, fa_s1_c81_n347_c;
    logic fa_s1_c81_n348_s, fa_s1_c81_n348_c;
    logic fa_s1_c81_n349_s, fa_s1_c81_n349_c;
    logic fa_s1_c82_n350_s, fa_s1_c82_n350_c;
    logic fa_s1_c82_n351_s, fa_s1_c82_n351_c;
    logic fa_s1_c82_n352_s, fa_s1_c82_n352_c;
    logic fa_s1_c82_n353_s, fa_s1_c82_n353_c;
    logic fa_s1_c82_n354_s, fa_s1_c82_n354_c;
    logic fa_s1_c82_n355_s, fa_s1_c82_n355_c;
    logic fa_s1_c82_n356_s, fa_s1_c82_n356_c;
    logic fa_s1_c83_n357_s, fa_s1_c83_n357_c;
    logic fa_s1_c83_n358_s, fa_s1_c83_n358_c;
    logic fa_s1_c83_n359_s, fa_s1_c83_n359_c;
    logic fa_s1_c83_n360_s, fa_s1_c83_n360_c;
    logic fa_s1_c83_n361_s, fa_s1_c83_n361_c;
    logic fa_s1_c83_n362_s, fa_s1_c83_n362_c;
    logic fa_s1_c83_n363_s, fa_s1_c83_n363_c;
    logic fa_s1_c84_n364_s, fa_s1_c84_n364_c;
    logic fa_s1_c84_n365_s, fa_s1_c84_n365_c;
    logic fa_s1_c84_n366_s, fa_s1_c84_n366_c;
    logic fa_s1_c84_n367_s, fa_s1_c84_n367_c;
    logic fa_s1_c84_n368_s, fa_s1_c84_n368_c;
    logic fa_s1_c84_n369_s, fa_s1_c84_n369_c;
    logic fa_s1_c84_n370_s, fa_s1_c84_n370_c;
    logic fa_s1_c85_n371_s, fa_s1_c85_n371_c;
    logic fa_s1_c85_n372_s, fa_s1_c85_n372_c;
    logic fa_s1_c85_n373_s, fa_s1_c85_n373_c;
    logic fa_s1_c85_n374_s, fa_s1_c85_n374_c;
    logic fa_s1_c85_n375_s, fa_s1_c85_n375_c;
    logic fa_s1_c85_n376_s, fa_s1_c85_n376_c;
    logic fa_s1_c85_n377_s, fa_s1_c85_n377_c;
    logic fa_s1_c86_n378_s, fa_s1_c86_n378_c;
    logic fa_s1_c86_n379_s, fa_s1_c86_n379_c;
    logic fa_s1_c86_n380_s, fa_s1_c86_n380_c;
    logic fa_s1_c86_n381_s, fa_s1_c86_n381_c;
    logic fa_s1_c86_n382_s, fa_s1_c86_n382_c;
    logic fa_s1_c86_n383_s, fa_s1_c86_n383_c;
    logic fa_s1_c86_n384_s, fa_s1_c86_n384_c;
    logic fa_s1_c87_n385_s, fa_s1_c87_n385_c;
    logic fa_s1_c87_n386_s, fa_s1_c87_n386_c;
    logic fa_s1_c87_n387_s, fa_s1_c87_n387_c;
    logic fa_s1_c87_n388_s, fa_s1_c87_n388_c;
    logic fa_s1_c87_n389_s, fa_s1_c87_n389_c;
    logic fa_s1_c87_n390_s, fa_s1_c87_n390_c;
    logic fa_s1_c87_n391_s, fa_s1_c87_n391_c;
    logic fa_s1_c88_n392_s, fa_s1_c88_n392_c;
    logic fa_s1_c88_n393_s, fa_s1_c88_n393_c;
    logic fa_s1_c88_n394_s, fa_s1_c88_n394_c;
    logic fa_s1_c88_n395_s, fa_s1_c88_n395_c;
    logic fa_s1_c88_n396_s, fa_s1_c88_n396_c;
    logic fa_s1_c88_n397_s, fa_s1_c88_n397_c;
    logic fa_s1_c88_n398_s, fa_s1_c88_n398_c;
    logic fa_s1_c89_n399_s, fa_s1_c89_n399_c;
    logic fa_s1_c89_n400_s, fa_s1_c89_n400_c;
    logic fa_s1_c89_n401_s, fa_s1_c89_n401_c;
    logic fa_s1_c89_n402_s, fa_s1_c89_n402_c;
    logic fa_s1_c89_n403_s, fa_s1_c89_n403_c;
    logic fa_s1_c89_n404_s, fa_s1_c89_n404_c;
    logic fa_s1_c89_n405_s, fa_s1_c89_n405_c;
    logic fa_s1_c90_n406_s, fa_s1_c90_n406_c;
    logic fa_s1_c90_n407_s, fa_s1_c90_n407_c;
    logic fa_s1_c90_n408_s, fa_s1_c90_n408_c;
    logic fa_s1_c90_n409_s, fa_s1_c90_n409_c;
    logic fa_s1_c90_n410_s, fa_s1_c90_n410_c;
    logic fa_s1_c90_n411_s, fa_s1_c90_n411_c;
    logic fa_s1_c90_n412_s, fa_s1_c90_n412_c;
    logic fa_s1_c91_n413_s, fa_s1_c91_n413_c;
    logic fa_s1_c91_n414_s, fa_s1_c91_n414_c;
    logic fa_s1_c91_n415_s, fa_s1_c91_n415_c;
    logic fa_s1_c91_n416_s, fa_s1_c91_n416_c;
    logic fa_s1_c91_n417_s, fa_s1_c91_n417_c;
    logic fa_s1_c91_n418_s, fa_s1_c91_n418_c;
    logic fa_s1_c91_n419_s, fa_s1_c91_n419_c;
    logic fa_s1_c92_n420_s, fa_s1_c92_n420_c;
    logic fa_s1_c92_n421_s, fa_s1_c92_n421_c;
    logic fa_s1_c92_n422_s, fa_s1_c92_n422_c;
    logic fa_s1_c92_n423_s, fa_s1_c92_n423_c;
    logic fa_s1_c92_n424_s, fa_s1_c92_n424_c;
    logic fa_s1_c92_n425_s, fa_s1_c92_n425_c;
    logic fa_s1_c92_n426_s, fa_s1_c92_n426_c;
    logic fa_s1_c93_n427_s, fa_s1_c93_n427_c;
    logic fa_s1_c93_n428_s, fa_s1_c93_n428_c;
    logic fa_s1_c93_n429_s, fa_s1_c93_n429_c;
    logic fa_s1_c93_n430_s, fa_s1_c93_n430_c;
    logic fa_s1_c93_n431_s, fa_s1_c93_n431_c;
    logic fa_s1_c93_n432_s, fa_s1_c93_n432_c;
    logic fa_s1_c93_n433_s, fa_s1_c93_n433_c;
    logic fa_s1_c94_n434_s, fa_s1_c94_n434_c;
    logic fa_s1_c94_n435_s, fa_s1_c94_n435_c;
    logic fa_s1_c94_n436_s, fa_s1_c94_n436_c;
    logic fa_s1_c94_n437_s, fa_s1_c94_n437_c;
    logic fa_s1_c94_n438_s, fa_s1_c94_n438_c;
    logic fa_s1_c94_n439_s, fa_s1_c94_n439_c;
    logic fa_s1_c94_n440_s, fa_s1_c94_n440_c;
    logic fa_s1_c95_n441_s, fa_s1_c95_n441_c;
    logic fa_s1_c95_n442_s, fa_s1_c95_n442_c;
    logic fa_s1_c95_n443_s, fa_s1_c95_n443_c;
    logic fa_s1_c95_n444_s, fa_s1_c95_n444_c;
    logic fa_s1_c95_n445_s, fa_s1_c95_n445_c;
    logic fa_s1_c95_n446_s, fa_s1_c95_n446_c;
    logic fa_s1_c95_n447_s, fa_s1_c95_n447_c;
    logic fa_s1_c96_n448_s, fa_s1_c96_n448_c;
    logic fa_s1_c96_n449_s, fa_s1_c96_n449_c;
    logic fa_s1_c96_n450_s, fa_s1_c96_n450_c;
    logic fa_s1_c96_n451_s, fa_s1_c96_n451_c;
    logic fa_s1_c96_n452_s, fa_s1_c96_n452_c;
    logic fa_s1_c96_n453_s, fa_s1_c96_n453_c;
    logic fa_s1_c96_n454_s, fa_s1_c96_n454_c;
    logic fa_s1_c97_n455_s, fa_s1_c97_n455_c;
    logic fa_s1_c97_n456_s, fa_s1_c97_n456_c;
    logic fa_s1_c97_n457_s, fa_s1_c97_n457_c;
    logic fa_s1_c97_n458_s, fa_s1_c97_n458_c;
    logic fa_s1_c97_n459_s, fa_s1_c97_n459_c;
    logic fa_s1_c97_n460_s, fa_s1_c97_n460_c;
    logic fa_s1_c97_n461_s, fa_s1_c97_n461_c;
    logic fa_s1_c98_n462_s, fa_s1_c98_n462_c;
    logic fa_s1_c98_n463_s, fa_s1_c98_n463_c;
    logic fa_s1_c98_n464_s, fa_s1_c98_n464_c;
    logic fa_s1_c98_n465_s, fa_s1_c98_n465_c;
    logic fa_s1_c98_n466_s, fa_s1_c98_n466_c;
    logic fa_s1_c98_n467_s, fa_s1_c98_n467_c;
    logic fa_s1_c98_n468_s, fa_s1_c98_n468_c;
    logic fa_s1_c99_n469_s, fa_s1_c99_n469_c;
    logic fa_s1_c99_n470_s, fa_s1_c99_n470_c;
    logic fa_s1_c99_n471_s, fa_s1_c99_n471_c;
    logic fa_s1_c99_n472_s, fa_s1_c99_n472_c;
    logic fa_s1_c99_n473_s, fa_s1_c99_n473_c;
    logic fa_s1_c99_n474_s, fa_s1_c99_n474_c;
    logic fa_s1_c99_n475_s, fa_s1_c99_n475_c;
    logic fa_s1_c100_n476_s, fa_s1_c100_n476_c;
    logic fa_s1_c100_n477_s, fa_s1_c100_n477_c;
    logic fa_s1_c100_n478_s, fa_s1_c100_n478_c;
    logic fa_s1_c100_n479_s, fa_s1_c100_n479_c;
    logic fa_s1_c100_n480_s, fa_s1_c100_n480_c;
    logic fa_s1_c100_n481_s, fa_s1_c100_n481_c;
    logic fa_s1_c100_n482_s, fa_s1_c100_n482_c;
    logic fa_s1_c101_n483_s, fa_s1_c101_n483_c;
    logic fa_s1_c101_n484_s, fa_s1_c101_n484_c;
    logic fa_s1_c101_n485_s, fa_s1_c101_n485_c;
    logic fa_s1_c101_n486_s, fa_s1_c101_n486_c;
    logic fa_s1_c101_n487_s, fa_s1_c101_n487_c;
    logic fa_s1_c101_n488_s, fa_s1_c101_n488_c;
    logic fa_s1_c101_n489_s, fa_s1_c101_n489_c;
    logic fa_s1_c102_n490_s, fa_s1_c102_n490_c;
    logic fa_s1_c102_n491_s, fa_s1_c102_n491_c;
    logic fa_s1_c102_n492_s, fa_s1_c102_n492_c;
    logic fa_s1_c102_n493_s, fa_s1_c102_n493_c;
    logic fa_s1_c102_n494_s, fa_s1_c102_n494_c;
    logic fa_s1_c102_n495_s, fa_s1_c102_n495_c;
    logic fa_s1_c102_n496_s, fa_s1_c102_n496_c;
    logic fa_s1_c103_n497_s, fa_s1_c103_n497_c;
    logic fa_s1_c103_n498_s, fa_s1_c103_n498_c;
    logic fa_s1_c103_n499_s, fa_s1_c103_n499_c;
    logic fa_s1_c103_n500_s, fa_s1_c103_n500_c;
    logic fa_s1_c103_n501_s, fa_s1_c103_n501_c;
    logic fa_s1_c103_n502_s, fa_s1_c103_n502_c;
    logic fa_s1_c103_n503_s, fa_s1_c103_n503_c;
    logic fa_s1_c104_n504_s, fa_s1_c104_n504_c;
    logic fa_s1_c104_n505_s, fa_s1_c104_n505_c;
    logic fa_s1_c104_n506_s, fa_s1_c104_n506_c;
    logic fa_s1_c104_n507_s, fa_s1_c104_n507_c;
    logic fa_s1_c104_n508_s, fa_s1_c104_n508_c;
    logic fa_s1_c104_n509_s, fa_s1_c104_n509_c;
    logic fa_s1_c104_n510_s, fa_s1_c104_n510_c;
    logic fa_s1_c105_n511_s, fa_s1_c105_n511_c;
    logic fa_s1_c105_n512_s, fa_s1_c105_n512_c;
    logic fa_s1_c105_n513_s, fa_s1_c105_n513_c;
    logic fa_s1_c105_n514_s, fa_s1_c105_n514_c;
    logic fa_s1_c105_n515_s, fa_s1_c105_n515_c;
    logic fa_s1_c105_n516_s, fa_s1_c105_n516_c;
    logic fa_s1_c105_n517_s, fa_s1_c105_n517_c;
    logic fa_s1_c106_n518_s, fa_s1_c106_n518_c;
    logic fa_s1_c106_n519_s, fa_s1_c106_n519_c;
    logic fa_s1_c106_n520_s, fa_s1_c106_n520_c;
    logic fa_s1_c106_n521_s, fa_s1_c106_n521_c;
    logic fa_s1_c106_n522_s, fa_s1_c106_n522_c;
    logic fa_s1_c106_n523_s, fa_s1_c106_n523_c;
    logic fa_s1_c106_n524_s, fa_s1_c106_n524_c;
    logic fa_s1_c107_n525_s, fa_s1_c107_n525_c;
    logic fa_s1_c107_n526_s, fa_s1_c107_n526_c;
    logic fa_s1_c107_n527_s, fa_s1_c107_n527_c;
    logic fa_s1_c107_n528_s, fa_s1_c107_n528_c;
    logic fa_s1_c107_n529_s, fa_s1_c107_n529_c;
    logic fa_s1_c107_n530_s, fa_s1_c107_n530_c;
    logic fa_s1_c107_n531_s, fa_s1_c107_n531_c;
    logic fa_s1_c108_n532_s, fa_s1_c108_n532_c;
    logic fa_s1_c108_n533_s, fa_s1_c108_n533_c;
    logic fa_s1_c108_n534_s, fa_s1_c108_n534_c;
    logic fa_s1_c108_n535_s, fa_s1_c108_n535_c;
    logic fa_s1_c108_n536_s, fa_s1_c108_n536_c;
    logic fa_s1_c108_n537_s, fa_s1_c108_n537_c;
    logic fa_s1_c108_n538_s, fa_s1_c108_n538_c;
    logic fa_s1_c109_n539_s, fa_s1_c109_n539_c;
    logic fa_s1_c109_n540_s, fa_s1_c109_n540_c;
    logic fa_s1_c109_n541_s, fa_s1_c109_n541_c;
    logic fa_s1_c109_n542_s, fa_s1_c109_n542_c;
    logic fa_s1_c109_n543_s, fa_s1_c109_n543_c;
    logic fa_s1_c109_n544_s, fa_s1_c109_n544_c;
    logic fa_s1_c109_n545_s, fa_s1_c109_n545_c;
    logic fa_s1_c110_n546_s, fa_s1_c110_n546_c;
    logic fa_s1_c110_n547_s, fa_s1_c110_n547_c;
    logic fa_s1_c110_n548_s, fa_s1_c110_n548_c;
    logic fa_s1_c110_n549_s, fa_s1_c110_n549_c;
    logic fa_s1_c110_n550_s, fa_s1_c110_n550_c;
    logic fa_s1_c110_n551_s, fa_s1_c110_n551_c;
    logic fa_s1_c110_n552_s, fa_s1_c110_n552_c;
    logic fa_s1_c111_n553_s, fa_s1_c111_n553_c;
    logic fa_s1_c111_n554_s, fa_s1_c111_n554_c;
    logic fa_s1_c111_n555_s, fa_s1_c111_n555_c;
    logic fa_s1_c111_n556_s, fa_s1_c111_n556_c;
    logic fa_s1_c111_n557_s, fa_s1_c111_n557_c;
    logic fa_s1_c111_n558_s, fa_s1_c111_n558_c;
    logic fa_s1_c111_n559_s, fa_s1_c111_n559_c;
    logic fa_s1_c112_n560_s, fa_s1_c112_n560_c;
    logic fa_s1_c112_n561_s, fa_s1_c112_n561_c;
    logic fa_s1_c112_n562_s, fa_s1_c112_n562_c;
    logic fa_s1_c112_n563_s, fa_s1_c112_n563_c;
    logic fa_s1_c112_n564_s, fa_s1_c112_n564_c;
    logic fa_s1_c112_n565_s, fa_s1_c112_n565_c;
    logic fa_s1_c112_n566_s, fa_s1_c112_n566_c;
    logic fa_s1_c113_n567_s, fa_s1_c113_n567_c;
    logic fa_s1_c113_n568_s, fa_s1_c113_n568_c;
    logic fa_s1_c113_n569_s, fa_s1_c113_n569_c;
    logic fa_s1_c113_n570_s, fa_s1_c113_n570_c;
    logic fa_s1_c113_n571_s, fa_s1_c113_n571_c;
    logic fa_s1_c113_n572_s, fa_s1_c113_n572_c;
    logic fa_s1_c113_n573_s, fa_s1_c113_n573_c;
    logic fa_s1_c114_n574_s, fa_s1_c114_n574_c;
    logic fa_s1_c114_n575_s, fa_s1_c114_n575_c;
    logic fa_s1_c114_n576_s, fa_s1_c114_n576_c;
    logic fa_s1_c114_n577_s, fa_s1_c114_n577_c;
    logic fa_s1_c114_n578_s, fa_s1_c114_n578_c;
    logic fa_s1_c114_n579_s, fa_s1_c114_n579_c;
    logic fa_s1_c114_n580_s, fa_s1_c114_n580_c;
    logic fa_s1_c115_n581_s, fa_s1_c115_n581_c;
    logic fa_s1_c115_n582_s, fa_s1_c115_n582_c;
    logic fa_s1_c115_n583_s, fa_s1_c115_n583_c;
    logic fa_s1_c115_n584_s, fa_s1_c115_n584_c;
    logic fa_s1_c115_n585_s, fa_s1_c115_n585_c;
    logic fa_s1_c115_n586_s, fa_s1_c115_n586_c;
    logic fa_s1_c115_n587_s, fa_s1_c115_n587_c;
    logic fa_s1_c116_n588_s, fa_s1_c116_n588_c;
    logic fa_s1_c116_n589_s, fa_s1_c116_n589_c;
    logic fa_s1_c116_n590_s, fa_s1_c116_n590_c;
    logic fa_s1_c116_n591_s, fa_s1_c116_n591_c;
    logic fa_s1_c116_n592_s, fa_s1_c116_n592_c;
    logic fa_s1_c116_n593_s, fa_s1_c116_n593_c;
    logic fa_s1_c116_n594_s, fa_s1_c116_n594_c;
    logic fa_s1_c117_n595_s, fa_s1_c117_n595_c;
    logic fa_s1_c117_n596_s, fa_s1_c117_n596_c;
    logic fa_s1_c117_n597_s, fa_s1_c117_n597_c;
    logic fa_s1_c117_n598_s, fa_s1_c117_n598_c;
    logic fa_s1_c117_n599_s, fa_s1_c117_n599_c;
    logic fa_s1_c117_n600_s, fa_s1_c117_n600_c;
    logic fa_s1_c117_n601_s, fa_s1_c117_n601_c;
    logic fa_s1_c118_n602_s, fa_s1_c118_n602_c;
    logic fa_s1_c118_n603_s, fa_s1_c118_n603_c;
    logic fa_s1_c118_n604_s, fa_s1_c118_n604_c;
    logic fa_s1_c118_n605_s, fa_s1_c118_n605_c;
    logic fa_s1_c118_n606_s, fa_s1_c118_n606_c;
    logic fa_s1_c118_n607_s, fa_s1_c118_n607_c;
    logic fa_s1_c118_n608_s, fa_s1_c118_n608_c;
    logic fa_s1_c119_n609_s, fa_s1_c119_n609_c;
    logic fa_s1_c119_n610_s, fa_s1_c119_n610_c;
    logic fa_s1_c119_n611_s, fa_s1_c119_n611_c;
    logic fa_s1_c119_n612_s, fa_s1_c119_n612_c;
    logic fa_s1_c119_n613_s, fa_s1_c119_n613_c;
    logic fa_s1_c119_n614_s, fa_s1_c119_n614_c;
    logic fa_s1_c119_n615_s, fa_s1_c119_n615_c;
    logic fa_s1_c120_n616_s, fa_s1_c120_n616_c;
    logic fa_s1_c120_n617_s, fa_s1_c120_n617_c;
    logic fa_s1_c120_n618_s, fa_s1_c120_n618_c;
    logic fa_s1_c120_n619_s, fa_s1_c120_n619_c;
    logic fa_s1_c120_n620_s, fa_s1_c120_n620_c;
    logic fa_s1_c120_n621_s, fa_s1_c120_n621_c;
    logic fa_s1_c120_n622_s, fa_s1_c120_n622_c;
    logic fa_s1_c121_n623_s, fa_s1_c121_n623_c;
    logic fa_s1_c121_n624_s, fa_s1_c121_n624_c;
    logic fa_s1_c121_n625_s, fa_s1_c121_n625_c;
    logic fa_s1_c121_n626_s, fa_s1_c121_n626_c;
    logic fa_s1_c121_n627_s, fa_s1_c121_n627_c;
    logic fa_s1_c121_n628_s, fa_s1_c121_n628_c;
    logic fa_s1_c121_n629_s, fa_s1_c121_n629_c;
    logic fa_s1_c122_n630_s, fa_s1_c122_n630_c;
    logic fa_s1_c122_n631_s, fa_s1_c122_n631_c;
    logic fa_s1_c122_n632_s, fa_s1_c122_n632_c;
    logic fa_s1_c122_n633_s, fa_s1_c122_n633_c;
    logic fa_s1_c122_n634_s, fa_s1_c122_n634_c;
    logic fa_s1_c122_n635_s, fa_s1_c122_n635_c;
    logic fa_s1_c122_n636_s, fa_s1_c122_n636_c;
    logic fa_s1_c123_n637_s, fa_s1_c123_n637_c;
    logic fa_s1_c123_n638_s, fa_s1_c123_n638_c;
    logic fa_s1_c123_n639_s, fa_s1_c123_n639_c;
    logic fa_s1_c123_n640_s, fa_s1_c123_n640_c;
    logic fa_s1_c123_n641_s, fa_s1_c123_n641_c;
    logic fa_s1_c123_n642_s, fa_s1_c123_n642_c;
    logic fa_s1_c123_n643_s, fa_s1_c123_n643_c;
    logic fa_s1_c124_n644_s, fa_s1_c124_n644_c;
    logic fa_s1_c124_n645_s, fa_s1_c124_n645_c;
    logic fa_s1_c124_n646_s, fa_s1_c124_n646_c;
    logic fa_s1_c124_n647_s, fa_s1_c124_n647_c;
    logic fa_s1_c124_n648_s, fa_s1_c124_n648_c;
    logic fa_s1_c124_n649_s, fa_s1_c124_n649_c;
    logic fa_s1_c124_n650_s, fa_s1_c124_n650_c;
    logic fa_s1_c125_n651_s, fa_s1_c125_n651_c;
    logic fa_s1_c125_n652_s, fa_s1_c125_n652_c;
    logic fa_s1_c125_n653_s, fa_s1_c125_n653_c;
    logic fa_s1_c125_n654_s, fa_s1_c125_n654_c;
    logic fa_s1_c125_n655_s, fa_s1_c125_n655_c;
    logic fa_s1_c125_n656_s, fa_s1_c125_n656_c;
    logic fa_s1_c125_n657_s, fa_s1_c125_n657_c;
    logic fa_s1_c126_n658_s, fa_s1_c126_n658_c;
    logic fa_s1_c126_n659_s, fa_s1_c126_n659_c;
    logic fa_s1_c126_n660_s, fa_s1_c126_n660_c;
    logic fa_s1_c126_n661_s, fa_s1_c126_n661_c;
    logic fa_s1_c126_n662_s, fa_s1_c126_n662_c;
    logic fa_s1_c126_n663_s, fa_s1_c126_n663_c;
    logic fa_s1_c126_n664_s, fa_s1_c126_n664_c;
    logic fa_s2_c4_n0_s, fa_s2_c4_n0_c;
    logic fa_s2_c9_n1_s, fa_s2_c9_n1_c;
    logic fa_s2_c10_n2_s, fa_s2_c10_n2_c;
    logic fa_s2_c11_n3_s, fa_s2_c11_n3_c;
    logic fa_s2_c12_n4_s, fa_s2_c12_n4_c;
    logic fa_s2_c13_n5_s, fa_s2_c13_n5_c;
    logic fa_s2_c14_n6_s, fa_s2_c14_n6_c;
    logic fa_s2_c15_n7_s, fa_s2_c15_n7_c;
    logic fa_s2_c16_n8_s, fa_s2_c16_n8_c;
    logic fa_s2_c17_n9_s, fa_s2_c17_n9_c;
    logic fa_s2_c18_n10_s, fa_s2_c18_n10_c;
    logic fa_s2_c18_n11_s, fa_s2_c18_n11_c;
    logic fa_s2_c19_n12_s, fa_s2_c19_n12_c;
    logic fa_s2_c20_n13_s, fa_s2_c20_n13_c;
    logic fa_s2_c21_n14_s, fa_s2_c21_n14_c;
    logic fa_s2_c22_n15_s, fa_s2_c22_n15_c;
    logic fa_s2_c22_n16_s, fa_s2_c22_n16_c;
    logic fa_s2_c23_n17_s, fa_s2_c23_n17_c;
    logic fa_s2_c23_n18_s, fa_s2_c23_n18_c;
    logic fa_s2_c24_n19_s, fa_s2_c24_n19_c;
    logic fa_s2_c24_n20_s, fa_s2_c24_n20_c;
    logic fa_s2_c25_n21_s, fa_s2_c25_n21_c;
    logic fa_s2_c25_n22_s, fa_s2_c25_n22_c;
    logic fa_s2_c26_n23_s, fa_s2_c26_n23_c;
    logic fa_s2_c26_n24_s, fa_s2_c26_n24_c;
    logic fa_s2_c27_n25_s, fa_s2_c27_n25_c;
    logic fa_s2_c27_n26_s, fa_s2_c27_n26_c;
    logic fa_s2_c28_n27_s, fa_s2_c28_n27_c;
    logic fa_s2_c28_n28_s, fa_s2_c28_n28_c;
    logic fa_s2_c29_n29_s, fa_s2_c29_n29_c;
    logic fa_s2_c29_n30_s, fa_s2_c29_n30_c;
    logic fa_s2_c30_n31_s, fa_s2_c30_n31_c;
    logic fa_s2_c30_n32_s, fa_s2_c30_n32_c;
    logic fa_s2_c31_n33_s, fa_s2_c31_n33_c;
    logic fa_s2_c31_n34_s, fa_s2_c31_n34_c;
    logic fa_s2_c31_n35_s, fa_s2_c31_n35_c;
    logic fa_s2_c32_n36_s, fa_s2_c32_n36_c;
    logic fa_s2_c32_n37_s, fa_s2_c32_n37_c;
    logic fa_s2_c33_n38_s, fa_s2_c33_n38_c;
    logic fa_s2_c33_n39_s, fa_s2_c33_n39_c;
    logic fa_s2_c34_n40_s, fa_s2_c34_n40_c;
    logic fa_s2_c34_n41_s, fa_s2_c34_n41_c;
    logic fa_s2_c35_n42_s, fa_s2_c35_n42_c;
    logic fa_s2_c35_n43_s, fa_s2_c35_n43_c;
    logic fa_s2_c36_n44_s, fa_s2_c36_n44_c;
    logic fa_s2_c36_n45_s, fa_s2_c36_n45_c;
    logic fa_s2_c36_n46_s, fa_s2_c36_n46_c;
    logic fa_s2_c37_n47_s, fa_s2_c37_n47_c;
    logic fa_s2_c37_n48_s, fa_s2_c37_n48_c;
    logic fa_s2_c37_n49_s, fa_s2_c37_n49_c;
    logic fa_s2_c38_n50_s, fa_s2_c38_n50_c;
    logic fa_s2_c38_n51_s, fa_s2_c38_n51_c;
    logic fa_s2_c38_n52_s, fa_s2_c38_n52_c;
    logic fa_s2_c39_n53_s, fa_s2_c39_n53_c;
    logic fa_s2_c39_n54_s, fa_s2_c39_n54_c;
    logic fa_s2_c39_n55_s, fa_s2_c39_n55_c;
    logic fa_s2_c40_n56_s, fa_s2_c40_n56_c;
    logic fa_s2_c40_n57_s, fa_s2_c40_n57_c;
    logic fa_s2_c40_n58_s, fa_s2_c40_n58_c;
    logic fa_s2_c41_n59_s, fa_s2_c41_n59_c;
    logic fa_s2_c41_n60_s, fa_s2_c41_n60_c;
    logic fa_s2_c41_n61_s, fa_s2_c41_n61_c;
    logic fa_s2_c42_n62_s, fa_s2_c42_n62_c;
    logic fa_s2_c42_n63_s, fa_s2_c42_n63_c;
    logic fa_s2_c42_n64_s, fa_s2_c42_n64_c;
    logic fa_s2_c43_n65_s, fa_s2_c43_n65_c;
    logic fa_s2_c43_n66_s, fa_s2_c43_n66_c;
    logic fa_s2_c43_n67_s, fa_s2_c43_n67_c;
    logic fa_s2_c44_n68_s, fa_s2_c44_n68_c;
    logic fa_s2_c44_n69_s, fa_s2_c44_n69_c;
    logic fa_s2_c44_n70_s, fa_s2_c44_n70_c;
    logic fa_s2_c45_n71_s, fa_s2_c45_n71_c;
    logic fa_s2_c45_n72_s, fa_s2_c45_n72_c;
    logic fa_s2_c45_n73_s, fa_s2_c45_n73_c;
    logic fa_s2_c45_n74_s, fa_s2_c45_n74_c;
    logic fa_s2_c46_n75_s, fa_s2_c46_n75_c;
    logic fa_s2_c46_n76_s, fa_s2_c46_n76_c;
    logic fa_s2_c46_n77_s, fa_s2_c46_n77_c;
    logic fa_s2_c47_n78_s, fa_s2_c47_n78_c;
    logic fa_s2_c47_n79_s, fa_s2_c47_n79_c;
    logic fa_s2_c47_n80_s, fa_s2_c47_n80_c;
    logic fa_s2_c48_n81_s, fa_s2_c48_n81_c;
    logic fa_s2_c48_n82_s, fa_s2_c48_n82_c;
    logic fa_s2_c48_n83_s, fa_s2_c48_n83_c;
    logic fa_s2_c49_n84_s, fa_s2_c49_n84_c;
    logic fa_s2_c49_n85_s, fa_s2_c49_n85_c;
    logic fa_s2_c49_n86_s, fa_s2_c49_n86_c;
    logic fa_s2_c49_n87_s, fa_s2_c49_n87_c;
    logic fa_s2_c50_n88_s, fa_s2_c50_n88_c;
    logic fa_s2_c50_n89_s, fa_s2_c50_n89_c;
    logic fa_s2_c50_n90_s, fa_s2_c50_n90_c;
    logic fa_s2_c50_n91_s, fa_s2_c50_n91_c;
    logic fa_s2_c51_n92_s, fa_s2_c51_n92_c;
    logic fa_s2_c51_n93_s, fa_s2_c51_n93_c;
    logic fa_s2_c51_n94_s, fa_s2_c51_n94_c;
    logic fa_s2_c51_n95_s, fa_s2_c51_n95_c;
    logic fa_s2_c52_n96_s, fa_s2_c52_n96_c;
    logic fa_s2_c52_n97_s, fa_s2_c52_n97_c;
    logic fa_s2_c52_n98_s, fa_s2_c52_n98_c;
    logic fa_s2_c52_n99_s, fa_s2_c52_n99_c;
    logic fa_s2_c53_n100_s, fa_s2_c53_n100_c;
    logic fa_s2_c53_n101_s, fa_s2_c53_n101_c;
    logic fa_s2_c53_n102_s, fa_s2_c53_n102_c;
    logic fa_s2_c53_n103_s, fa_s2_c53_n103_c;
    logic fa_s2_c54_n104_s, fa_s2_c54_n104_c;
    logic fa_s2_c54_n105_s, fa_s2_c54_n105_c;
    logic fa_s2_c54_n106_s, fa_s2_c54_n106_c;
    logic fa_s2_c54_n107_s, fa_s2_c54_n107_c;
    logic fa_s2_c55_n108_s, fa_s2_c55_n108_c;
    logic fa_s2_c55_n109_s, fa_s2_c55_n109_c;
    logic fa_s2_c55_n110_s, fa_s2_c55_n110_c;
    logic fa_s2_c55_n111_s, fa_s2_c55_n111_c;
    logic fa_s2_c56_n112_s, fa_s2_c56_n112_c;
    logic fa_s2_c56_n113_s, fa_s2_c56_n113_c;
    logic fa_s2_c56_n114_s, fa_s2_c56_n114_c;
    logic fa_s2_c56_n115_s, fa_s2_c56_n115_c;
    logic fa_s2_c57_n116_s, fa_s2_c57_n116_c;
    logic fa_s2_c57_n117_s, fa_s2_c57_n117_c;
    logic fa_s2_c57_n118_s, fa_s2_c57_n118_c;
    logic fa_s2_c57_n119_s, fa_s2_c57_n119_c;
    logic fa_s2_c58_n120_s, fa_s2_c58_n120_c;
    logic fa_s2_c58_n121_s, fa_s2_c58_n121_c;
    logic fa_s2_c58_n122_s, fa_s2_c58_n122_c;
    logic fa_s2_c58_n123_s, fa_s2_c58_n123_c;
    logic fa_s2_c58_n124_s, fa_s2_c58_n124_c;
    logic fa_s2_c59_n125_s, fa_s2_c59_n125_c;
    logic fa_s2_c59_n126_s, fa_s2_c59_n126_c;
    logic fa_s2_c59_n127_s, fa_s2_c59_n127_c;
    logic fa_s2_c59_n128_s, fa_s2_c59_n128_c;
    logic fa_s2_c60_n129_s, fa_s2_c60_n129_c;
    logic fa_s2_c60_n130_s, fa_s2_c60_n130_c;
    logic fa_s2_c60_n131_s, fa_s2_c60_n131_c;
    logic fa_s2_c60_n132_s, fa_s2_c60_n132_c;
    logic fa_s2_c61_n133_s, fa_s2_c61_n133_c;
    logic fa_s2_c61_n134_s, fa_s2_c61_n134_c;
    logic fa_s2_c61_n135_s, fa_s2_c61_n135_c;
    logic fa_s2_c61_n136_s, fa_s2_c61_n136_c;
    logic fa_s2_c62_n137_s, fa_s2_c62_n137_c;
    logic fa_s2_c62_n138_s, fa_s2_c62_n138_c;
    logic fa_s2_c62_n139_s, fa_s2_c62_n139_c;
    logic fa_s2_c62_n140_s, fa_s2_c62_n140_c;
    logic fa_s2_c63_n141_s, fa_s2_c63_n141_c;
    logic fa_s2_c63_n142_s, fa_s2_c63_n142_c;
    logic fa_s2_c63_n143_s, fa_s2_c63_n143_c;
    logic fa_s2_c63_n144_s, fa_s2_c63_n144_c;
    logic fa_s2_c63_n145_s, fa_s2_c63_n145_c;
    logic fa_s2_c64_n146_s, fa_s2_c64_n146_c;
    logic fa_s2_c64_n147_s, fa_s2_c64_n147_c;
    logic fa_s2_c64_n148_s, fa_s2_c64_n148_c;
    logic fa_s2_c64_n149_s, fa_s2_c64_n149_c;
    logic fa_s2_c65_n150_s, fa_s2_c65_n150_c;
    logic fa_s2_c65_n151_s, fa_s2_c65_n151_c;
    logic fa_s2_c65_n152_s, fa_s2_c65_n152_c;
    logic fa_s2_c65_n153_s, fa_s2_c65_n153_c;
    logic fa_s2_c65_n154_s, fa_s2_c65_n154_c;
    logic fa_s2_c66_n155_s, fa_s2_c66_n155_c;
    logic fa_s2_c66_n156_s, fa_s2_c66_n156_c;
    logic fa_s2_c66_n157_s, fa_s2_c66_n157_c;
    logic fa_s2_c66_n158_s, fa_s2_c66_n158_c;
    logic fa_s2_c67_n159_s, fa_s2_c67_n159_c;
    logic fa_s2_c67_n160_s, fa_s2_c67_n160_c;
    logic fa_s2_c67_n161_s, fa_s2_c67_n161_c;
    logic fa_s2_c67_n162_s, fa_s2_c67_n162_c;
    logic fa_s2_c67_n163_s, fa_s2_c67_n163_c;
    logic fa_s2_c68_n164_s, fa_s2_c68_n164_c;
    logic fa_s2_c68_n165_s, fa_s2_c68_n165_c;
    logic fa_s2_c68_n166_s, fa_s2_c68_n166_c;
    logic fa_s2_c68_n167_s, fa_s2_c68_n167_c;
    logic fa_s2_c69_n168_s, fa_s2_c69_n168_c;
    logic fa_s2_c69_n169_s, fa_s2_c69_n169_c;
    logic fa_s2_c69_n170_s, fa_s2_c69_n170_c;
    logic fa_s2_c69_n171_s, fa_s2_c69_n171_c;
    logic fa_s2_c69_n172_s, fa_s2_c69_n172_c;
    logic fa_s2_c70_n173_s, fa_s2_c70_n173_c;
    logic fa_s2_c70_n174_s, fa_s2_c70_n174_c;
    logic fa_s2_c70_n175_s, fa_s2_c70_n175_c;
    logic fa_s2_c70_n176_s, fa_s2_c70_n176_c;
    logic fa_s2_c71_n177_s, fa_s2_c71_n177_c;
    logic fa_s2_c71_n178_s, fa_s2_c71_n178_c;
    logic fa_s2_c71_n179_s, fa_s2_c71_n179_c;
    logic fa_s2_c71_n180_s, fa_s2_c71_n180_c;
    logic fa_s2_c71_n181_s, fa_s2_c71_n181_c;
    logic fa_s2_c72_n182_s, fa_s2_c72_n182_c;
    logic fa_s2_c72_n183_s, fa_s2_c72_n183_c;
    logic fa_s2_c72_n184_s, fa_s2_c72_n184_c;
    logic fa_s2_c72_n185_s, fa_s2_c72_n185_c;
    logic fa_s2_c73_n186_s, fa_s2_c73_n186_c;
    logic fa_s2_c73_n187_s, fa_s2_c73_n187_c;
    logic fa_s2_c73_n188_s, fa_s2_c73_n188_c;
    logic fa_s2_c73_n189_s, fa_s2_c73_n189_c;
    logic fa_s2_c73_n190_s, fa_s2_c73_n190_c;
    logic fa_s2_c74_n191_s, fa_s2_c74_n191_c;
    logic fa_s2_c74_n192_s, fa_s2_c74_n192_c;
    logic fa_s2_c74_n193_s, fa_s2_c74_n193_c;
    logic fa_s2_c74_n194_s, fa_s2_c74_n194_c;
    logic fa_s2_c75_n195_s, fa_s2_c75_n195_c;
    logic fa_s2_c75_n196_s, fa_s2_c75_n196_c;
    logic fa_s2_c75_n197_s, fa_s2_c75_n197_c;
    logic fa_s2_c75_n198_s, fa_s2_c75_n198_c;
    logic fa_s2_c75_n199_s, fa_s2_c75_n199_c;
    logic fa_s2_c76_n200_s, fa_s2_c76_n200_c;
    logic fa_s2_c76_n201_s, fa_s2_c76_n201_c;
    logic fa_s2_c76_n202_s, fa_s2_c76_n202_c;
    logic fa_s2_c76_n203_s, fa_s2_c76_n203_c;
    logic fa_s2_c77_n204_s, fa_s2_c77_n204_c;
    logic fa_s2_c77_n205_s, fa_s2_c77_n205_c;
    logic fa_s2_c77_n206_s, fa_s2_c77_n206_c;
    logic fa_s2_c77_n207_s, fa_s2_c77_n207_c;
    logic fa_s2_c77_n208_s, fa_s2_c77_n208_c;
    logic fa_s2_c78_n209_s, fa_s2_c78_n209_c;
    logic fa_s2_c78_n210_s, fa_s2_c78_n210_c;
    logic fa_s2_c78_n211_s, fa_s2_c78_n211_c;
    logic fa_s2_c78_n212_s, fa_s2_c78_n212_c;
    logic fa_s2_c79_n213_s, fa_s2_c79_n213_c;
    logic fa_s2_c79_n214_s, fa_s2_c79_n214_c;
    logic fa_s2_c79_n215_s, fa_s2_c79_n215_c;
    logic fa_s2_c79_n216_s, fa_s2_c79_n216_c;
    logic fa_s2_c79_n217_s, fa_s2_c79_n217_c;
    logic fa_s2_c80_n218_s, fa_s2_c80_n218_c;
    logic fa_s2_c80_n219_s, fa_s2_c80_n219_c;
    logic fa_s2_c80_n220_s, fa_s2_c80_n220_c;
    logic fa_s2_c80_n221_s, fa_s2_c80_n221_c;
    logic fa_s2_c81_n222_s, fa_s2_c81_n222_c;
    logic fa_s2_c81_n223_s, fa_s2_c81_n223_c;
    logic fa_s2_c81_n224_s, fa_s2_c81_n224_c;
    logic fa_s2_c81_n225_s, fa_s2_c81_n225_c;
    logic fa_s2_c81_n226_s, fa_s2_c81_n226_c;
    logic fa_s2_c82_n227_s, fa_s2_c82_n227_c;
    logic fa_s2_c82_n228_s, fa_s2_c82_n228_c;
    logic fa_s2_c82_n229_s, fa_s2_c82_n229_c;
    logic fa_s2_c82_n230_s, fa_s2_c82_n230_c;
    logic fa_s2_c83_n231_s, fa_s2_c83_n231_c;
    logic fa_s2_c83_n232_s, fa_s2_c83_n232_c;
    logic fa_s2_c83_n233_s, fa_s2_c83_n233_c;
    logic fa_s2_c83_n234_s, fa_s2_c83_n234_c;
    logic fa_s2_c83_n235_s, fa_s2_c83_n235_c;
    logic fa_s2_c84_n236_s, fa_s2_c84_n236_c;
    logic fa_s2_c84_n237_s, fa_s2_c84_n237_c;
    logic fa_s2_c84_n238_s, fa_s2_c84_n238_c;
    logic fa_s2_c84_n239_s, fa_s2_c84_n239_c;
    logic fa_s2_c85_n240_s, fa_s2_c85_n240_c;
    logic fa_s2_c85_n241_s, fa_s2_c85_n241_c;
    logic fa_s2_c85_n242_s, fa_s2_c85_n242_c;
    logic fa_s2_c85_n243_s, fa_s2_c85_n243_c;
    logic fa_s2_c85_n244_s, fa_s2_c85_n244_c;
    logic fa_s2_c86_n245_s, fa_s2_c86_n245_c;
    logic fa_s2_c86_n246_s, fa_s2_c86_n246_c;
    logic fa_s2_c86_n247_s, fa_s2_c86_n247_c;
    logic fa_s2_c86_n248_s, fa_s2_c86_n248_c;
    logic fa_s2_c87_n249_s, fa_s2_c87_n249_c;
    logic fa_s2_c87_n250_s, fa_s2_c87_n250_c;
    logic fa_s2_c87_n251_s, fa_s2_c87_n251_c;
    logic fa_s2_c87_n252_s, fa_s2_c87_n252_c;
    logic fa_s2_c87_n253_s, fa_s2_c87_n253_c;
    logic fa_s2_c88_n254_s, fa_s2_c88_n254_c;
    logic fa_s2_c88_n255_s, fa_s2_c88_n255_c;
    logic fa_s2_c88_n256_s, fa_s2_c88_n256_c;
    logic fa_s2_c88_n257_s, fa_s2_c88_n257_c;
    logic fa_s2_c89_n258_s, fa_s2_c89_n258_c;
    logic fa_s2_c89_n259_s, fa_s2_c89_n259_c;
    logic fa_s2_c89_n260_s, fa_s2_c89_n260_c;
    logic fa_s2_c89_n261_s, fa_s2_c89_n261_c;
    logic fa_s2_c89_n262_s, fa_s2_c89_n262_c;
    logic fa_s2_c90_n263_s, fa_s2_c90_n263_c;
    logic fa_s2_c90_n264_s, fa_s2_c90_n264_c;
    logic fa_s2_c90_n265_s, fa_s2_c90_n265_c;
    logic fa_s2_c90_n266_s, fa_s2_c90_n266_c;
    logic fa_s2_c91_n267_s, fa_s2_c91_n267_c;
    logic fa_s2_c91_n268_s, fa_s2_c91_n268_c;
    logic fa_s2_c91_n269_s, fa_s2_c91_n269_c;
    logic fa_s2_c91_n270_s, fa_s2_c91_n270_c;
    logic fa_s2_c91_n271_s, fa_s2_c91_n271_c;
    logic fa_s2_c92_n272_s, fa_s2_c92_n272_c;
    logic fa_s2_c92_n273_s, fa_s2_c92_n273_c;
    logic fa_s2_c92_n274_s, fa_s2_c92_n274_c;
    logic fa_s2_c92_n275_s, fa_s2_c92_n275_c;
    logic fa_s2_c93_n276_s, fa_s2_c93_n276_c;
    logic fa_s2_c93_n277_s, fa_s2_c93_n277_c;
    logic fa_s2_c93_n278_s, fa_s2_c93_n278_c;
    logic fa_s2_c93_n279_s, fa_s2_c93_n279_c;
    logic fa_s2_c93_n280_s, fa_s2_c93_n280_c;
    logic fa_s2_c94_n281_s, fa_s2_c94_n281_c;
    logic fa_s2_c94_n282_s, fa_s2_c94_n282_c;
    logic fa_s2_c94_n283_s, fa_s2_c94_n283_c;
    logic fa_s2_c94_n284_s, fa_s2_c94_n284_c;
    logic fa_s2_c95_n285_s, fa_s2_c95_n285_c;
    logic fa_s2_c95_n286_s, fa_s2_c95_n286_c;
    logic fa_s2_c95_n287_s, fa_s2_c95_n287_c;
    logic fa_s2_c95_n288_s, fa_s2_c95_n288_c;
    logic fa_s2_c95_n289_s, fa_s2_c95_n289_c;
    logic fa_s2_c96_n290_s, fa_s2_c96_n290_c;
    logic fa_s2_c96_n291_s, fa_s2_c96_n291_c;
    logic fa_s2_c96_n292_s, fa_s2_c96_n292_c;
    logic fa_s2_c96_n293_s, fa_s2_c96_n293_c;
    logic fa_s2_c97_n294_s, fa_s2_c97_n294_c;
    logic fa_s2_c97_n295_s, fa_s2_c97_n295_c;
    logic fa_s2_c97_n296_s, fa_s2_c97_n296_c;
    logic fa_s2_c97_n297_s, fa_s2_c97_n297_c;
    logic fa_s2_c97_n298_s, fa_s2_c97_n298_c;
    logic fa_s2_c98_n299_s, fa_s2_c98_n299_c;
    logic fa_s2_c98_n300_s, fa_s2_c98_n300_c;
    logic fa_s2_c98_n301_s, fa_s2_c98_n301_c;
    logic fa_s2_c98_n302_s, fa_s2_c98_n302_c;
    logic fa_s2_c99_n303_s, fa_s2_c99_n303_c;
    logic fa_s2_c99_n304_s, fa_s2_c99_n304_c;
    logic fa_s2_c99_n305_s, fa_s2_c99_n305_c;
    logic fa_s2_c99_n306_s, fa_s2_c99_n306_c;
    logic fa_s2_c99_n307_s, fa_s2_c99_n307_c;
    logic fa_s2_c100_n308_s, fa_s2_c100_n308_c;
    logic fa_s2_c100_n309_s, fa_s2_c100_n309_c;
    logic fa_s2_c100_n310_s, fa_s2_c100_n310_c;
    logic fa_s2_c100_n311_s, fa_s2_c100_n311_c;
    logic fa_s2_c101_n312_s, fa_s2_c101_n312_c;
    logic fa_s2_c101_n313_s, fa_s2_c101_n313_c;
    logic fa_s2_c101_n314_s, fa_s2_c101_n314_c;
    logic fa_s2_c101_n315_s, fa_s2_c101_n315_c;
    logic fa_s2_c101_n316_s, fa_s2_c101_n316_c;
    logic fa_s2_c102_n317_s, fa_s2_c102_n317_c;
    logic fa_s2_c102_n318_s, fa_s2_c102_n318_c;
    logic fa_s2_c102_n319_s, fa_s2_c102_n319_c;
    logic fa_s2_c102_n320_s, fa_s2_c102_n320_c;
    logic fa_s2_c103_n321_s, fa_s2_c103_n321_c;
    logic fa_s2_c103_n322_s, fa_s2_c103_n322_c;
    logic fa_s2_c103_n323_s, fa_s2_c103_n323_c;
    logic fa_s2_c103_n324_s, fa_s2_c103_n324_c;
    logic fa_s2_c103_n325_s, fa_s2_c103_n325_c;
    logic fa_s2_c104_n326_s, fa_s2_c104_n326_c;
    logic fa_s2_c104_n327_s, fa_s2_c104_n327_c;
    logic fa_s2_c104_n328_s, fa_s2_c104_n328_c;
    logic fa_s2_c104_n329_s, fa_s2_c104_n329_c;
    logic fa_s2_c105_n330_s, fa_s2_c105_n330_c;
    logic fa_s2_c105_n331_s, fa_s2_c105_n331_c;
    logic fa_s2_c105_n332_s, fa_s2_c105_n332_c;
    logic fa_s2_c105_n333_s, fa_s2_c105_n333_c;
    logic fa_s2_c105_n334_s, fa_s2_c105_n334_c;
    logic fa_s2_c106_n335_s, fa_s2_c106_n335_c;
    logic fa_s2_c106_n336_s, fa_s2_c106_n336_c;
    logic fa_s2_c106_n337_s, fa_s2_c106_n337_c;
    logic fa_s2_c106_n338_s, fa_s2_c106_n338_c;
    logic fa_s2_c107_n339_s, fa_s2_c107_n339_c;
    logic fa_s2_c107_n340_s, fa_s2_c107_n340_c;
    logic fa_s2_c107_n341_s, fa_s2_c107_n341_c;
    logic fa_s2_c107_n342_s, fa_s2_c107_n342_c;
    logic fa_s2_c107_n343_s, fa_s2_c107_n343_c;
    logic fa_s2_c108_n344_s, fa_s2_c108_n344_c;
    logic fa_s2_c108_n345_s, fa_s2_c108_n345_c;
    logic fa_s2_c108_n346_s, fa_s2_c108_n346_c;
    logic fa_s2_c108_n347_s, fa_s2_c108_n347_c;
    logic fa_s2_c109_n348_s, fa_s2_c109_n348_c;
    logic fa_s2_c109_n349_s, fa_s2_c109_n349_c;
    logic fa_s2_c109_n350_s, fa_s2_c109_n350_c;
    logic fa_s2_c109_n351_s, fa_s2_c109_n351_c;
    logic fa_s2_c109_n352_s, fa_s2_c109_n352_c;
    logic fa_s2_c110_n353_s, fa_s2_c110_n353_c;
    logic fa_s2_c110_n354_s, fa_s2_c110_n354_c;
    logic fa_s2_c110_n355_s, fa_s2_c110_n355_c;
    logic fa_s2_c110_n356_s, fa_s2_c110_n356_c;
    logic fa_s2_c111_n357_s, fa_s2_c111_n357_c;
    logic fa_s2_c111_n358_s, fa_s2_c111_n358_c;
    logic fa_s2_c111_n359_s, fa_s2_c111_n359_c;
    logic fa_s2_c111_n360_s, fa_s2_c111_n360_c;
    logic fa_s2_c111_n361_s, fa_s2_c111_n361_c;
    logic fa_s2_c112_n362_s, fa_s2_c112_n362_c;
    logic fa_s2_c112_n363_s, fa_s2_c112_n363_c;
    logic fa_s2_c112_n364_s, fa_s2_c112_n364_c;
    logic fa_s2_c112_n365_s, fa_s2_c112_n365_c;
    logic fa_s2_c113_n366_s, fa_s2_c113_n366_c;
    logic fa_s2_c113_n367_s, fa_s2_c113_n367_c;
    logic fa_s2_c113_n368_s, fa_s2_c113_n368_c;
    logic fa_s2_c113_n369_s, fa_s2_c113_n369_c;
    logic fa_s2_c113_n370_s, fa_s2_c113_n370_c;
    logic fa_s2_c114_n371_s, fa_s2_c114_n371_c;
    logic fa_s2_c114_n372_s, fa_s2_c114_n372_c;
    logic fa_s2_c114_n373_s, fa_s2_c114_n373_c;
    logic fa_s2_c114_n374_s, fa_s2_c114_n374_c;
    logic fa_s2_c115_n375_s, fa_s2_c115_n375_c;
    logic fa_s2_c115_n376_s, fa_s2_c115_n376_c;
    logic fa_s2_c115_n377_s, fa_s2_c115_n377_c;
    logic fa_s2_c115_n378_s, fa_s2_c115_n378_c;
    logic fa_s2_c115_n379_s, fa_s2_c115_n379_c;
    logic fa_s2_c116_n380_s, fa_s2_c116_n380_c;
    logic fa_s2_c116_n381_s, fa_s2_c116_n381_c;
    logic fa_s2_c116_n382_s, fa_s2_c116_n382_c;
    logic fa_s2_c116_n383_s, fa_s2_c116_n383_c;
    logic fa_s2_c117_n384_s, fa_s2_c117_n384_c;
    logic fa_s2_c117_n385_s, fa_s2_c117_n385_c;
    logic fa_s2_c117_n386_s, fa_s2_c117_n386_c;
    logic fa_s2_c117_n387_s, fa_s2_c117_n387_c;
    logic fa_s2_c117_n388_s, fa_s2_c117_n388_c;
    logic fa_s2_c118_n389_s, fa_s2_c118_n389_c;
    logic fa_s2_c118_n390_s, fa_s2_c118_n390_c;
    logic fa_s2_c118_n391_s, fa_s2_c118_n391_c;
    logic fa_s2_c118_n392_s, fa_s2_c118_n392_c;
    logic fa_s2_c119_n393_s, fa_s2_c119_n393_c;
    logic fa_s2_c119_n394_s, fa_s2_c119_n394_c;
    logic fa_s2_c119_n395_s, fa_s2_c119_n395_c;
    logic fa_s2_c119_n396_s, fa_s2_c119_n396_c;
    logic fa_s2_c119_n397_s, fa_s2_c119_n397_c;
    logic fa_s2_c120_n398_s, fa_s2_c120_n398_c;
    logic fa_s2_c120_n399_s, fa_s2_c120_n399_c;
    logic fa_s2_c120_n400_s, fa_s2_c120_n400_c;
    logic fa_s2_c120_n401_s, fa_s2_c120_n401_c;
    logic fa_s2_c121_n402_s, fa_s2_c121_n402_c;
    logic fa_s2_c121_n403_s, fa_s2_c121_n403_c;
    logic fa_s2_c121_n404_s, fa_s2_c121_n404_c;
    logic fa_s2_c121_n405_s, fa_s2_c121_n405_c;
    logic fa_s2_c121_n406_s, fa_s2_c121_n406_c;
    logic fa_s2_c122_n407_s, fa_s2_c122_n407_c;
    logic fa_s2_c122_n408_s, fa_s2_c122_n408_c;
    logic fa_s2_c122_n409_s, fa_s2_c122_n409_c;
    logic fa_s2_c122_n410_s, fa_s2_c122_n410_c;
    logic fa_s2_c123_n411_s, fa_s2_c123_n411_c;
    logic fa_s2_c123_n412_s, fa_s2_c123_n412_c;
    logic fa_s2_c123_n413_s, fa_s2_c123_n413_c;
    logic fa_s2_c123_n414_s, fa_s2_c123_n414_c;
    logic fa_s2_c123_n415_s, fa_s2_c123_n415_c;
    logic fa_s2_c124_n416_s, fa_s2_c124_n416_c;
    logic fa_s2_c124_n417_s, fa_s2_c124_n417_c;
    logic fa_s2_c124_n418_s, fa_s2_c124_n418_c;
    logic fa_s2_c124_n419_s, fa_s2_c124_n419_c;
    logic fa_s2_c125_n420_s, fa_s2_c125_n420_c;
    logic fa_s2_c125_n421_s, fa_s2_c125_n421_c;
    logic fa_s2_c125_n422_s, fa_s2_c125_n422_c;
    logic fa_s2_c125_n423_s, fa_s2_c125_n423_c;
    logic fa_s2_c125_n424_s, fa_s2_c125_n424_c;
    logic fa_s2_c126_n425_s, fa_s2_c126_n425_c;
    logic fa_s2_c126_n426_s, fa_s2_c126_n426_c;
    logic fa_s2_c126_n427_s, fa_s2_c126_n427_c;
    logic fa_s2_c126_n428_s, fa_s2_c126_n428_c;
    logic fa_s3_c5_n0_s, fa_s3_c5_n0_c;
    logic fa_s3_c13_n1_s, fa_s3_c13_n1_c;
    logic fa_s3_c14_n2_s, fa_s3_c14_n2_c;
    logic fa_s3_c15_n3_s, fa_s3_c15_n3_c;
    logic fa_s3_c16_n4_s, fa_s3_c16_n4_c;
    logic fa_s3_c17_n5_s, fa_s3_c17_n5_c;
    logic fa_s3_c18_n6_s, fa_s3_c18_n6_c;
    logic fa_s3_c19_n7_s, fa_s3_c19_n7_c;
    logic fa_s3_c20_n8_s, fa_s3_c20_n8_c;
    logic fa_s3_c21_n9_s, fa_s3_c21_n9_c;
    logic fa_s3_c22_n10_s, fa_s3_c22_n10_c;
    logic fa_s3_c23_n11_s, fa_s3_c23_n11_c;
    logic fa_s3_c24_n12_s, fa_s3_c24_n12_c;
    logic fa_s3_c25_n13_s, fa_s3_c25_n13_c;
    logic fa_s3_c26_n14_s, fa_s3_c26_n14_c;
    logic fa_s3_c27_n15_s, fa_s3_c27_n15_c;
    logic fa_s3_c27_n16_s, fa_s3_c27_n16_c;
    logic fa_s3_c28_n17_s, fa_s3_c28_n17_c;
    logic fa_s3_c29_n18_s, fa_s3_c29_n18_c;
    logic fa_s3_c30_n19_s, fa_s3_c30_n19_c;
    logic fa_s3_c31_n20_s, fa_s3_c31_n20_c;
    logic fa_s3_c32_n21_s, fa_s3_c32_n21_c;
    logic fa_s3_c32_n22_s, fa_s3_c32_n22_c;
    logic fa_s3_c33_n23_s, fa_s3_c33_n23_c;
    logic fa_s3_c33_n24_s, fa_s3_c33_n24_c;
    logic fa_s3_c34_n25_s, fa_s3_c34_n25_c;
    logic fa_s3_c34_n26_s, fa_s3_c34_n26_c;
    logic fa_s3_c35_n27_s, fa_s3_c35_n27_c;
    logic fa_s3_c35_n28_s, fa_s3_c35_n28_c;
    logic fa_s3_c36_n29_s, fa_s3_c36_n29_c;
    logic fa_s3_c36_n30_s, fa_s3_c36_n30_c;
    logic fa_s3_c37_n31_s, fa_s3_c37_n31_c;
    logic fa_s3_c37_n32_s, fa_s3_c37_n32_c;
    logic fa_s3_c38_n33_s, fa_s3_c38_n33_c;
    logic fa_s3_c38_n34_s, fa_s3_c38_n34_c;
    logic fa_s3_c39_n35_s, fa_s3_c39_n35_c;
    logic fa_s3_c39_n36_s, fa_s3_c39_n36_c;
    logic fa_s3_c40_n37_s, fa_s3_c40_n37_c;
    logic fa_s3_c40_n38_s, fa_s3_c40_n38_c;
    logic fa_s3_c41_n39_s, fa_s3_c41_n39_c;
    logic fa_s3_c41_n40_s, fa_s3_c41_n40_c;
    logic fa_s3_c42_n41_s, fa_s3_c42_n41_c;
    logic fa_s3_c42_n42_s, fa_s3_c42_n42_c;
    logic fa_s3_c43_n43_s, fa_s3_c43_n43_c;
    logic fa_s3_c43_n44_s, fa_s3_c43_n44_c;
    logic fa_s3_c44_n45_s, fa_s3_c44_n45_c;
    logic fa_s3_c44_n46_s, fa_s3_c44_n46_c;
    logic fa_s3_c45_n47_s, fa_s3_c45_n47_c;
    logic fa_s3_c45_n48_s, fa_s3_c45_n48_c;
    logic fa_s3_c46_n49_s, fa_s3_c46_n49_c;
    logic fa_s3_c46_n50_s, fa_s3_c46_n50_c;
    logic fa_s3_c46_n51_s, fa_s3_c46_n51_c;
    logic fa_s3_c47_n52_s, fa_s3_c47_n52_c;
    logic fa_s3_c47_n53_s, fa_s3_c47_n53_c;
    logic fa_s3_c48_n54_s, fa_s3_c48_n54_c;
    logic fa_s3_c48_n55_s, fa_s3_c48_n55_c;
    logic fa_s3_c49_n56_s, fa_s3_c49_n56_c;
    logic fa_s3_c49_n57_s, fa_s3_c49_n57_c;
    logic fa_s3_c50_n58_s, fa_s3_c50_n58_c;
    logic fa_s3_c50_n59_s, fa_s3_c50_n59_c;
    logic fa_s3_c51_n60_s, fa_s3_c51_n60_c;
    logic fa_s3_c51_n61_s, fa_s3_c51_n61_c;
    logic fa_s3_c52_n62_s, fa_s3_c52_n62_c;
    logic fa_s3_c52_n63_s, fa_s3_c52_n63_c;
    logic fa_s3_c53_n64_s, fa_s3_c53_n64_c;
    logic fa_s3_c53_n65_s, fa_s3_c53_n65_c;
    logic fa_s3_c54_n66_s, fa_s3_c54_n66_c;
    logic fa_s3_c54_n67_s, fa_s3_c54_n67_c;
    logic fa_s3_c54_n68_s, fa_s3_c54_n68_c;
    logic fa_s3_c55_n69_s, fa_s3_c55_n69_c;
    logic fa_s3_c55_n70_s, fa_s3_c55_n70_c;
    logic fa_s3_c55_n71_s, fa_s3_c55_n71_c;
    logic fa_s3_c56_n72_s, fa_s3_c56_n72_c;
    logic fa_s3_c56_n73_s, fa_s3_c56_n73_c;
    logic fa_s3_c56_n74_s, fa_s3_c56_n74_c;
    logic fa_s3_c57_n75_s, fa_s3_c57_n75_c;
    logic fa_s3_c57_n76_s, fa_s3_c57_n76_c;
    logic fa_s3_c57_n77_s, fa_s3_c57_n77_c;
    logic fa_s3_c58_n78_s, fa_s3_c58_n78_c;
    logic fa_s3_c58_n79_s, fa_s3_c58_n79_c;
    logic fa_s3_c58_n80_s, fa_s3_c58_n80_c;
    logic fa_s3_c59_n81_s, fa_s3_c59_n81_c;
    logic fa_s3_c59_n82_s, fa_s3_c59_n82_c;
    logic fa_s3_c59_n83_s, fa_s3_c59_n83_c;
    logic fa_s3_c60_n84_s, fa_s3_c60_n84_c;
    logic fa_s3_c60_n85_s, fa_s3_c60_n85_c;
    logic fa_s3_c60_n86_s, fa_s3_c60_n86_c;
    logic fa_s3_c61_n87_s, fa_s3_c61_n87_c;
    logic fa_s3_c61_n88_s, fa_s3_c61_n88_c;
    logic fa_s3_c61_n89_s, fa_s3_c61_n89_c;
    logic fa_s3_c62_n90_s, fa_s3_c62_n90_c;
    logic fa_s3_c62_n91_s, fa_s3_c62_n91_c;
    logic fa_s3_c62_n92_s, fa_s3_c62_n92_c;
    logic fa_s3_c63_n93_s, fa_s3_c63_n93_c;
    logic fa_s3_c63_n94_s, fa_s3_c63_n94_c;
    logic fa_s3_c63_n95_s, fa_s3_c63_n95_c;
    logic fa_s3_c64_n96_s, fa_s3_c64_n96_c;
    logic fa_s3_c64_n97_s, fa_s3_c64_n97_c;
    logic fa_s3_c64_n98_s, fa_s3_c64_n98_c;
    logic fa_s3_c65_n99_s, fa_s3_c65_n99_c;
    logic fa_s3_c65_n100_s, fa_s3_c65_n100_c;
    logic fa_s3_c65_n101_s, fa_s3_c65_n101_c;
    logic fa_s3_c66_n102_s, fa_s3_c66_n102_c;
    logic fa_s3_c66_n103_s, fa_s3_c66_n103_c;
    logic fa_s3_c66_n104_s, fa_s3_c66_n104_c;
    logic fa_s3_c67_n105_s, fa_s3_c67_n105_c;
    logic fa_s3_c67_n106_s, fa_s3_c67_n106_c;
    logic fa_s3_c67_n107_s, fa_s3_c67_n107_c;
    logic fa_s3_c68_n108_s, fa_s3_c68_n108_c;
    logic fa_s3_c68_n109_s, fa_s3_c68_n109_c;
    logic fa_s3_c68_n110_s, fa_s3_c68_n110_c;
    logic fa_s3_c69_n111_s, fa_s3_c69_n111_c;
    logic fa_s3_c69_n112_s, fa_s3_c69_n112_c;
    logic fa_s3_c69_n113_s, fa_s3_c69_n113_c;
    logic fa_s3_c70_n114_s, fa_s3_c70_n114_c;
    logic fa_s3_c70_n115_s, fa_s3_c70_n115_c;
    logic fa_s3_c70_n116_s, fa_s3_c70_n116_c;
    logic fa_s3_c71_n117_s, fa_s3_c71_n117_c;
    logic fa_s3_c71_n118_s, fa_s3_c71_n118_c;
    logic fa_s3_c71_n119_s, fa_s3_c71_n119_c;
    logic fa_s3_c72_n120_s, fa_s3_c72_n120_c;
    logic fa_s3_c72_n121_s, fa_s3_c72_n121_c;
    logic fa_s3_c72_n122_s, fa_s3_c72_n122_c;
    logic fa_s3_c73_n123_s, fa_s3_c73_n123_c;
    logic fa_s3_c73_n124_s, fa_s3_c73_n124_c;
    logic fa_s3_c73_n125_s, fa_s3_c73_n125_c;
    logic fa_s3_c74_n126_s, fa_s3_c74_n126_c;
    logic fa_s3_c74_n127_s, fa_s3_c74_n127_c;
    logic fa_s3_c74_n128_s, fa_s3_c74_n128_c;
    logic fa_s3_c75_n129_s, fa_s3_c75_n129_c;
    logic fa_s3_c75_n130_s, fa_s3_c75_n130_c;
    logic fa_s3_c75_n131_s, fa_s3_c75_n131_c;
    logic fa_s3_c76_n132_s, fa_s3_c76_n132_c;
    logic fa_s3_c76_n133_s, fa_s3_c76_n133_c;
    logic fa_s3_c76_n134_s, fa_s3_c76_n134_c;
    logic fa_s3_c77_n135_s, fa_s3_c77_n135_c;
    logic fa_s3_c77_n136_s, fa_s3_c77_n136_c;
    logic fa_s3_c77_n137_s, fa_s3_c77_n137_c;
    logic fa_s3_c78_n138_s, fa_s3_c78_n138_c;
    logic fa_s3_c78_n139_s, fa_s3_c78_n139_c;
    logic fa_s3_c78_n140_s, fa_s3_c78_n140_c;
    logic fa_s3_c79_n141_s, fa_s3_c79_n141_c;
    logic fa_s3_c79_n142_s, fa_s3_c79_n142_c;
    logic fa_s3_c79_n143_s, fa_s3_c79_n143_c;
    logic fa_s3_c80_n144_s, fa_s3_c80_n144_c;
    logic fa_s3_c80_n145_s, fa_s3_c80_n145_c;
    logic fa_s3_c80_n146_s, fa_s3_c80_n146_c;
    logic fa_s3_c81_n147_s, fa_s3_c81_n147_c;
    logic fa_s3_c81_n148_s, fa_s3_c81_n148_c;
    logic fa_s3_c81_n149_s, fa_s3_c81_n149_c;
    logic fa_s3_c82_n150_s, fa_s3_c82_n150_c;
    logic fa_s3_c82_n151_s, fa_s3_c82_n151_c;
    logic fa_s3_c82_n152_s, fa_s3_c82_n152_c;
    logic fa_s3_c83_n153_s, fa_s3_c83_n153_c;
    logic fa_s3_c83_n154_s, fa_s3_c83_n154_c;
    logic fa_s3_c83_n155_s, fa_s3_c83_n155_c;
    logic fa_s3_c84_n156_s, fa_s3_c84_n156_c;
    logic fa_s3_c84_n157_s, fa_s3_c84_n157_c;
    logic fa_s3_c84_n158_s, fa_s3_c84_n158_c;
    logic fa_s3_c85_n159_s, fa_s3_c85_n159_c;
    logic fa_s3_c85_n160_s, fa_s3_c85_n160_c;
    logic fa_s3_c85_n161_s, fa_s3_c85_n161_c;
    logic fa_s3_c86_n162_s, fa_s3_c86_n162_c;
    logic fa_s3_c86_n163_s, fa_s3_c86_n163_c;
    logic fa_s3_c86_n164_s, fa_s3_c86_n164_c;
    logic fa_s3_c87_n165_s, fa_s3_c87_n165_c;
    logic fa_s3_c87_n166_s, fa_s3_c87_n166_c;
    logic fa_s3_c87_n167_s, fa_s3_c87_n167_c;
    logic fa_s3_c88_n168_s, fa_s3_c88_n168_c;
    logic fa_s3_c88_n169_s, fa_s3_c88_n169_c;
    logic fa_s3_c88_n170_s, fa_s3_c88_n170_c;
    logic fa_s3_c89_n171_s, fa_s3_c89_n171_c;
    logic fa_s3_c89_n172_s, fa_s3_c89_n172_c;
    logic fa_s3_c89_n173_s, fa_s3_c89_n173_c;
    logic fa_s3_c90_n174_s, fa_s3_c90_n174_c;
    logic fa_s3_c90_n175_s, fa_s3_c90_n175_c;
    logic fa_s3_c90_n176_s, fa_s3_c90_n176_c;
    logic fa_s3_c91_n177_s, fa_s3_c91_n177_c;
    logic fa_s3_c91_n178_s, fa_s3_c91_n178_c;
    logic fa_s3_c91_n179_s, fa_s3_c91_n179_c;
    logic fa_s3_c92_n180_s, fa_s3_c92_n180_c;
    logic fa_s3_c92_n181_s, fa_s3_c92_n181_c;
    logic fa_s3_c92_n182_s, fa_s3_c92_n182_c;
    logic fa_s3_c93_n183_s, fa_s3_c93_n183_c;
    logic fa_s3_c93_n184_s, fa_s3_c93_n184_c;
    logic fa_s3_c93_n185_s, fa_s3_c93_n185_c;
    logic fa_s3_c94_n186_s, fa_s3_c94_n186_c;
    logic fa_s3_c94_n187_s, fa_s3_c94_n187_c;
    logic fa_s3_c94_n188_s, fa_s3_c94_n188_c;
    logic fa_s3_c95_n189_s, fa_s3_c95_n189_c;
    logic fa_s3_c95_n190_s, fa_s3_c95_n190_c;
    logic fa_s3_c95_n191_s, fa_s3_c95_n191_c;
    logic fa_s3_c96_n192_s, fa_s3_c96_n192_c;
    logic fa_s3_c96_n193_s, fa_s3_c96_n193_c;
    logic fa_s3_c96_n194_s, fa_s3_c96_n194_c;
    logic fa_s3_c97_n195_s, fa_s3_c97_n195_c;
    logic fa_s3_c97_n196_s, fa_s3_c97_n196_c;
    logic fa_s3_c97_n197_s, fa_s3_c97_n197_c;
    logic fa_s3_c98_n198_s, fa_s3_c98_n198_c;
    logic fa_s3_c98_n199_s, fa_s3_c98_n199_c;
    logic fa_s3_c98_n200_s, fa_s3_c98_n200_c;
    logic fa_s3_c99_n201_s, fa_s3_c99_n201_c;
    logic fa_s3_c99_n202_s, fa_s3_c99_n202_c;
    logic fa_s3_c99_n203_s, fa_s3_c99_n203_c;
    logic fa_s3_c100_n204_s, fa_s3_c100_n204_c;
    logic fa_s3_c100_n205_s, fa_s3_c100_n205_c;
    logic fa_s3_c100_n206_s, fa_s3_c100_n206_c;
    logic fa_s3_c101_n207_s, fa_s3_c101_n207_c;
    logic fa_s3_c101_n208_s, fa_s3_c101_n208_c;
    logic fa_s3_c101_n209_s, fa_s3_c101_n209_c;
    logic fa_s3_c102_n210_s, fa_s3_c102_n210_c;
    logic fa_s3_c102_n211_s, fa_s3_c102_n211_c;
    logic fa_s3_c102_n212_s, fa_s3_c102_n212_c;
    logic fa_s3_c103_n213_s, fa_s3_c103_n213_c;
    logic fa_s3_c103_n214_s, fa_s3_c103_n214_c;
    logic fa_s3_c103_n215_s, fa_s3_c103_n215_c;
    logic fa_s3_c104_n216_s, fa_s3_c104_n216_c;
    logic fa_s3_c104_n217_s, fa_s3_c104_n217_c;
    logic fa_s3_c104_n218_s, fa_s3_c104_n218_c;
    logic fa_s3_c105_n219_s, fa_s3_c105_n219_c;
    logic fa_s3_c105_n220_s, fa_s3_c105_n220_c;
    logic fa_s3_c105_n221_s, fa_s3_c105_n221_c;
    logic fa_s3_c106_n222_s, fa_s3_c106_n222_c;
    logic fa_s3_c106_n223_s, fa_s3_c106_n223_c;
    logic fa_s3_c106_n224_s, fa_s3_c106_n224_c;
    logic fa_s3_c107_n225_s, fa_s3_c107_n225_c;
    logic fa_s3_c107_n226_s, fa_s3_c107_n226_c;
    logic fa_s3_c107_n227_s, fa_s3_c107_n227_c;
    logic fa_s3_c108_n228_s, fa_s3_c108_n228_c;
    logic fa_s3_c108_n229_s, fa_s3_c108_n229_c;
    logic fa_s3_c108_n230_s, fa_s3_c108_n230_c;
    logic fa_s3_c109_n231_s, fa_s3_c109_n231_c;
    logic fa_s3_c109_n232_s, fa_s3_c109_n232_c;
    logic fa_s3_c109_n233_s, fa_s3_c109_n233_c;
    logic fa_s3_c110_n234_s, fa_s3_c110_n234_c;
    logic fa_s3_c110_n235_s, fa_s3_c110_n235_c;
    logic fa_s3_c110_n236_s, fa_s3_c110_n236_c;
    logic fa_s3_c111_n237_s, fa_s3_c111_n237_c;
    logic fa_s3_c111_n238_s, fa_s3_c111_n238_c;
    logic fa_s3_c111_n239_s, fa_s3_c111_n239_c;
    logic fa_s3_c112_n240_s, fa_s3_c112_n240_c;
    logic fa_s3_c112_n241_s, fa_s3_c112_n241_c;
    logic fa_s3_c112_n242_s, fa_s3_c112_n242_c;
    logic fa_s3_c113_n243_s, fa_s3_c113_n243_c;
    logic fa_s3_c113_n244_s, fa_s3_c113_n244_c;
    logic fa_s3_c113_n245_s, fa_s3_c113_n245_c;
    logic fa_s3_c114_n246_s, fa_s3_c114_n246_c;
    logic fa_s3_c114_n247_s, fa_s3_c114_n247_c;
    logic fa_s3_c114_n248_s, fa_s3_c114_n248_c;
    logic fa_s3_c115_n249_s, fa_s3_c115_n249_c;
    logic fa_s3_c115_n250_s, fa_s3_c115_n250_c;
    logic fa_s3_c115_n251_s, fa_s3_c115_n251_c;
    logic fa_s3_c116_n252_s, fa_s3_c116_n252_c;
    logic fa_s3_c116_n253_s, fa_s3_c116_n253_c;
    logic fa_s3_c116_n254_s, fa_s3_c116_n254_c;
    logic fa_s3_c117_n255_s, fa_s3_c117_n255_c;
    logic fa_s3_c117_n256_s, fa_s3_c117_n256_c;
    logic fa_s3_c117_n257_s, fa_s3_c117_n257_c;
    logic fa_s3_c118_n258_s, fa_s3_c118_n258_c;
    logic fa_s3_c118_n259_s, fa_s3_c118_n259_c;
    logic fa_s3_c118_n260_s, fa_s3_c118_n260_c;
    logic fa_s3_c119_n261_s, fa_s3_c119_n261_c;
    logic fa_s3_c119_n262_s, fa_s3_c119_n262_c;
    logic fa_s3_c119_n263_s, fa_s3_c119_n263_c;
    logic fa_s3_c120_n264_s, fa_s3_c120_n264_c;
    logic fa_s3_c120_n265_s, fa_s3_c120_n265_c;
    logic fa_s3_c120_n266_s, fa_s3_c120_n266_c;
    logic fa_s3_c121_n267_s, fa_s3_c121_n267_c;
    logic fa_s3_c121_n268_s, fa_s3_c121_n268_c;
    logic fa_s3_c121_n269_s, fa_s3_c121_n269_c;
    logic fa_s3_c122_n270_s, fa_s3_c122_n270_c;
    logic fa_s3_c122_n271_s, fa_s3_c122_n271_c;
    logic fa_s3_c122_n272_s, fa_s3_c122_n272_c;
    logic fa_s3_c123_n273_s, fa_s3_c123_n273_c;
    logic fa_s3_c123_n274_s, fa_s3_c123_n274_c;
    logic fa_s3_c123_n275_s, fa_s3_c123_n275_c;
    logic fa_s3_c124_n276_s, fa_s3_c124_n276_c;
    logic fa_s3_c124_n277_s, fa_s3_c124_n277_c;
    logic fa_s3_c124_n278_s, fa_s3_c124_n278_c;
    logic fa_s3_c125_n279_s, fa_s3_c125_n279_c;
    logic fa_s3_c125_n280_s, fa_s3_c125_n280_c;
    logic fa_s3_c125_n281_s, fa_s3_c125_n281_c;
    logic fa_s3_c126_n282_s, fa_s3_c126_n282_c;
    logic fa_s3_c126_n283_s, fa_s3_c126_n283_c;
    logic fa_s3_c126_n284_s, fa_s3_c126_n284_c;
    logic fa_s4_c6_n0_s, fa_s4_c6_n0_c;
    logic fa_s4_c19_n1_s, fa_s4_c19_n1_c;
    logic fa_s4_c20_n2_s, fa_s4_c20_n2_c;
    logic fa_s4_c21_n3_s, fa_s4_c21_n3_c;
    logic fa_s4_c22_n4_s, fa_s4_c22_n4_c;
    logic fa_s4_c23_n5_s, fa_s4_c23_n5_c;
    logic fa_s4_c24_n6_s, fa_s4_c24_n6_c;
    logic fa_s4_c25_n7_s, fa_s4_c25_n7_c;
    logic fa_s4_c26_n8_s, fa_s4_c26_n8_c;
    logic fa_s4_c27_n9_s, fa_s4_c27_n9_c;
    logic fa_s4_c28_n10_s, fa_s4_c28_n10_c;
    logic fa_s4_c29_n11_s, fa_s4_c29_n11_c;
    logic fa_s4_c30_n12_s, fa_s4_c30_n12_c;
    logic fa_s4_c31_n13_s, fa_s4_c31_n13_c;
    logic fa_s4_c32_n14_s, fa_s4_c32_n14_c;
    logic fa_s4_c33_n15_s, fa_s4_c33_n15_c;
    logic fa_s4_c34_n16_s, fa_s4_c34_n16_c;
    logic fa_s4_c35_n17_s, fa_s4_c35_n17_c;
    logic fa_s4_c36_n18_s, fa_s4_c36_n18_c;
    logic fa_s4_c37_n19_s, fa_s4_c37_n19_c;
    logic fa_s4_c38_n20_s, fa_s4_c38_n20_c;
    logic fa_s4_c39_n21_s, fa_s4_c39_n21_c;
    logic fa_s4_c40_n22_s, fa_s4_c40_n22_c;
    logic fa_s4_c40_n23_s, fa_s4_c40_n23_c;
    logic fa_s4_c41_n24_s, fa_s4_c41_n24_c;
    logic fa_s4_c42_n25_s, fa_s4_c42_n25_c;
    logic fa_s4_c43_n26_s, fa_s4_c43_n26_c;
    logic fa_s4_c44_n27_s, fa_s4_c44_n27_c;
    logic fa_s4_c45_n28_s, fa_s4_c45_n28_c;
    logic fa_s4_c46_n29_s, fa_s4_c46_n29_c;
    logic fa_s4_c47_n30_s, fa_s4_c47_n30_c;
    logic fa_s4_c47_n31_s, fa_s4_c47_n31_c;
    logic fa_s4_c48_n32_s, fa_s4_c48_n32_c;
    logic fa_s4_c48_n33_s, fa_s4_c48_n33_c;
    logic fa_s4_c49_n34_s, fa_s4_c49_n34_c;
    logic fa_s4_c49_n35_s, fa_s4_c49_n35_c;
    logic fa_s4_c50_n36_s, fa_s4_c50_n36_c;
    logic fa_s4_c50_n37_s, fa_s4_c50_n37_c;
    logic fa_s4_c51_n38_s, fa_s4_c51_n38_c;
    logic fa_s4_c51_n39_s, fa_s4_c51_n39_c;
    logic fa_s4_c52_n40_s, fa_s4_c52_n40_c;
    logic fa_s4_c52_n41_s, fa_s4_c52_n41_c;
    logic fa_s4_c53_n42_s, fa_s4_c53_n42_c;
    logic fa_s4_c53_n43_s, fa_s4_c53_n43_c;
    logic fa_s4_c54_n44_s, fa_s4_c54_n44_c;
    logic fa_s4_c54_n45_s, fa_s4_c54_n45_c;
    logic fa_s4_c55_n46_s, fa_s4_c55_n46_c;
    logic fa_s4_c55_n47_s, fa_s4_c55_n47_c;
    logic fa_s4_c56_n48_s, fa_s4_c56_n48_c;
    logic fa_s4_c56_n49_s, fa_s4_c56_n49_c;
    logic fa_s4_c57_n50_s, fa_s4_c57_n50_c;
    logic fa_s4_c57_n51_s, fa_s4_c57_n51_c;
    logic fa_s4_c58_n52_s, fa_s4_c58_n52_c;
    logic fa_s4_c58_n53_s, fa_s4_c58_n53_c;
    logic fa_s4_c59_n54_s, fa_s4_c59_n54_c;
    logic fa_s4_c59_n55_s, fa_s4_c59_n55_c;
    logic fa_s4_c60_n56_s, fa_s4_c60_n56_c;
    logic fa_s4_c60_n57_s, fa_s4_c60_n57_c;
    logic fa_s4_c61_n58_s, fa_s4_c61_n58_c;
    logic fa_s4_c61_n59_s, fa_s4_c61_n59_c;
    logic fa_s4_c62_n60_s, fa_s4_c62_n60_c;
    logic fa_s4_c62_n61_s, fa_s4_c62_n61_c;
    logic fa_s4_c63_n62_s, fa_s4_c63_n62_c;
    logic fa_s4_c63_n63_s, fa_s4_c63_n63_c;
    logic fa_s4_c64_n64_s, fa_s4_c64_n64_c;
    logic fa_s4_c64_n65_s, fa_s4_c64_n65_c;
    logic fa_s4_c65_n66_s, fa_s4_c65_n66_c;
    logic fa_s4_c65_n67_s, fa_s4_c65_n67_c;
    logic fa_s4_c66_n68_s, fa_s4_c66_n68_c;
    logic fa_s4_c66_n69_s, fa_s4_c66_n69_c;
    logic fa_s4_c67_n70_s, fa_s4_c67_n70_c;
    logic fa_s4_c67_n71_s, fa_s4_c67_n71_c;
    logic fa_s4_c68_n72_s, fa_s4_c68_n72_c;
    logic fa_s4_c68_n73_s, fa_s4_c68_n73_c;
    logic fa_s4_c69_n74_s, fa_s4_c69_n74_c;
    logic fa_s4_c69_n75_s, fa_s4_c69_n75_c;
    logic fa_s4_c70_n76_s, fa_s4_c70_n76_c;
    logic fa_s4_c70_n77_s, fa_s4_c70_n77_c;
    logic fa_s4_c71_n78_s, fa_s4_c71_n78_c;
    logic fa_s4_c71_n79_s, fa_s4_c71_n79_c;
    logic fa_s4_c72_n80_s, fa_s4_c72_n80_c;
    logic fa_s4_c72_n81_s, fa_s4_c72_n81_c;
    logic fa_s4_c73_n82_s, fa_s4_c73_n82_c;
    logic fa_s4_c73_n83_s, fa_s4_c73_n83_c;
    logic fa_s4_c74_n84_s, fa_s4_c74_n84_c;
    logic fa_s4_c74_n85_s, fa_s4_c74_n85_c;
    logic fa_s4_c75_n86_s, fa_s4_c75_n86_c;
    logic fa_s4_c75_n87_s, fa_s4_c75_n87_c;
    logic fa_s4_c76_n88_s, fa_s4_c76_n88_c;
    logic fa_s4_c76_n89_s, fa_s4_c76_n89_c;
    logic fa_s4_c77_n90_s, fa_s4_c77_n90_c;
    logic fa_s4_c77_n91_s, fa_s4_c77_n91_c;
    logic fa_s4_c78_n92_s, fa_s4_c78_n92_c;
    logic fa_s4_c78_n93_s, fa_s4_c78_n93_c;
    logic fa_s4_c79_n94_s, fa_s4_c79_n94_c;
    logic fa_s4_c79_n95_s, fa_s4_c79_n95_c;
    logic fa_s4_c80_n96_s, fa_s4_c80_n96_c;
    logic fa_s4_c80_n97_s, fa_s4_c80_n97_c;
    logic fa_s4_c81_n98_s, fa_s4_c81_n98_c;
    logic fa_s4_c81_n99_s, fa_s4_c81_n99_c;
    logic fa_s4_c82_n100_s, fa_s4_c82_n100_c;
    logic fa_s4_c82_n101_s, fa_s4_c82_n101_c;
    logic fa_s4_c83_n102_s, fa_s4_c83_n102_c;
    logic fa_s4_c83_n103_s, fa_s4_c83_n103_c;
    logic fa_s4_c84_n104_s, fa_s4_c84_n104_c;
    logic fa_s4_c84_n105_s, fa_s4_c84_n105_c;
    logic fa_s4_c85_n106_s, fa_s4_c85_n106_c;
    logic fa_s4_c85_n107_s, fa_s4_c85_n107_c;
    logic fa_s4_c86_n108_s, fa_s4_c86_n108_c;
    logic fa_s4_c86_n109_s, fa_s4_c86_n109_c;
    logic fa_s4_c87_n110_s, fa_s4_c87_n110_c;
    logic fa_s4_c87_n111_s, fa_s4_c87_n111_c;
    logic fa_s4_c88_n112_s, fa_s4_c88_n112_c;
    logic fa_s4_c88_n113_s, fa_s4_c88_n113_c;
    logic fa_s4_c89_n114_s, fa_s4_c89_n114_c;
    logic fa_s4_c89_n115_s, fa_s4_c89_n115_c;
    logic fa_s4_c90_n116_s, fa_s4_c90_n116_c;
    logic fa_s4_c90_n117_s, fa_s4_c90_n117_c;
    logic fa_s4_c91_n118_s, fa_s4_c91_n118_c;
    logic fa_s4_c91_n119_s, fa_s4_c91_n119_c;
    logic fa_s4_c92_n120_s, fa_s4_c92_n120_c;
    logic fa_s4_c92_n121_s, fa_s4_c92_n121_c;
    logic fa_s4_c93_n122_s, fa_s4_c93_n122_c;
    logic fa_s4_c93_n123_s, fa_s4_c93_n123_c;
    logic fa_s4_c94_n124_s, fa_s4_c94_n124_c;
    logic fa_s4_c94_n125_s, fa_s4_c94_n125_c;
    logic fa_s4_c95_n126_s, fa_s4_c95_n126_c;
    logic fa_s4_c95_n127_s, fa_s4_c95_n127_c;
    logic fa_s4_c96_n128_s, fa_s4_c96_n128_c;
    logic fa_s4_c96_n129_s, fa_s4_c96_n129_c;
    logic fa_s4_c97_n130_s, fa_s4_c97_n130_c;
    logic fa_s4_c97_n131_s, fa_s4_c97_n131_c;
    logic fa_s4_c98_n132_s, fa_s4_c98_n132_c;
    logic fa_s4_c98_n133_s, fa_s4_c98_n133_c;
    logic fa_s4_c99_n134_s, fa_s4_c99_n134_c;
    logic fa_s4_c99_n135_s, fa_s4_c99_n135_c;
    logic fa_s4_c100_n136_s, fa_s4_c100_n136_c;
    logic fa_s4_c100_n137_s, fa_s4_c100_n137_c;
    logic fa_s4_c101_n138_s, fa_s4_c101_n138_c;
    logic fa_s4_c101_n139_s, fa_s4_c101_n139_c;
    logic fa_s4_c102_n140_s, fa_s4_c102_n140_c;
    logic fa_s4_c102_n141_s, fa_s4_c102_n141_c;
    logic fa_s4_c103_n142_s, fa_s4_c103_n142_c;
    logic fa_s4_c103_n143_s, fa_s4_c103_n143_c;
    logic fa_s4_c104_n144_s, fa_s4_c104_n144_c;
    logic fa_s4_c104_n145_s, fa_s4_c104_n145_c;
    logic fa_s4_c105_n146_s, fa_s4_c105_n146_c;
    logic fa_s4_c105_n147_s, fa_s4_c105_n147_c;
    logic fa_s4_c106_n148_s, fa_s4_c106_n148_c;
    logic fa_s4_c106_n149_s, fa_s4_c106_n149_c;
    logic fa_s4_c107_n150_s, fa_s4_c107_n150_c;
    logic fa_s4_c107_n151_s, fa_s4_c107_n151_c;
    logic fa_s4_c108_n152_s, fa_s4_c108_n152_c;
    logic fa_s4_c108_n153_s, fa_s4_c108_n153_c;
    logic fa_s4_c109_n154_s, fa_s4_c109_n154_c;
    logic fa_s4_c109_n155_s, fa_s4_c109_n155_c;
    logic fa_s4_c110_n156_s, fa_s4_c110_n156_c;
    logic fa_s4_c110_n157_s, fa_s4_c110_n157_c;
    logic fa_s4_c111_n158_s, fa_s4_c111_n158_c;
    logic fa_s4_c111_n159_s, fa_s4_c111_n159_c;
    logic fa_s4_c112_n160_s, fa_s4_c112_n160_c;
    logic fa_s4_c112_n161_s, fa_s4_c112_n161_c;
    logic fa_s4_c113_n162_s, fa_s4_c113_n162_c;
    logic fa_s4_c113_n163_s, fa_s4_c113_n163_c;
    logic fa_s4_c114_n164_s, fa_s4_c114_n164_c;
    logic fa_s4_c114_n165_s, fa_s4_c114_n165_c;
    logic fa_s4_c115_n166_s, fa_s4_c115_n166_c;
    logic fa_s4_c115_n167_s, fa_s4_c115_n167_c;
    logic fa_s4_c116_n168_s, fa_s4_c116_n168_c;
    logic fa_s4_c116_n169_s, fa_s4_c116_n169_c;
    logic fa_s4_c117_n170_s, fa_s4_c117_n170_c;
    logic fa_s4_c117_n171_s, fa_s4_c117_n171_c;
    logic fa_s4_c118_n172_s, fa_s4_c118_n172_c;
    logic fa_s4_c118_n173_s, fa_s4_c118_n173_c;
    logic fa_s4_c119_n174_s, fa_s4_c119_n174_c;
    logic fa_s4_c119_n175_s, fa_s4_c119_n175_c;
    logic fa_s4_c120_n176_s, fa_s4_c120_n176_c;
    logic fa_s4_c120_n177_s, fa_s4_c120_n177_c;
    logic fa_s4_c121_n178_s, fa_s4_c121_n178_c;
    logic fa_s4_c121_n179_s, fa_s4_c121_n179_c;
    logic fa_s4_c122_n180_s, fa_s4_c122_n180_c;
    logic fa_s4_c122_n181_s, fa_s4_c122_n181_c;
    logic fa_s4_c123_n182_s, fa_s4_c123_n182_c;
    logic fa_s4_c123_n183_s, fa_s4_c123_n183_c;
    logic fa_s4_c124_n184_s, fa_s4_c124_n184_c;
    logic fa_s4_c124_n185_s, fa_s4_c124_n185_c;
    logic fa_s4_c125_n186_s, fa_s4_c125_n186_c;
    logic fa_s4_c125_n187_s, fa_s4_c125_n187_c;
    logic fa_s4_c126_n188_s, fa_s4_c126_n188_c;
    logic fa_s4_c126_n189_s, fa_s4_c126_n189_c;
    logic fa_s5_c7_n0_s, fa_s5_c7_n0_c;
    logic fa_s5_c28_n1_s, fa_s5_c28_n1_c;
    logic fa_s5_c29_n2_s, fa_s5_c29_n2_c;
    logic fa_s5_c30_n3_s, fa_s5_c30_n3_c;
    logic fa_s5_c31_n4_s, fa_s5_c31_n4_c;
    logic fa_s5_c32_n5_s, fa_s5_c32_n5_c;
    logic fa_s5_c33_n6_s, fa_s5_c33_n6_c;
    logic fa_s5_c34_n7_s, fa_s5_c34_n7_c;
    logic fa_s5_c35_n8_s, fa_s5_c35_n8_c;
    logic fa_s5_c36_n9_s, fa_s5_c36_n9_c;
    logic fa_s5_c37_n10_s, fa_s5_c37_n10_c;
    logic fa_s5_c38_n11_s, fa_s5_c38_n11_c;
    logic fa_s5_c39_n12_s, fa_s5_c39_n12_c;
    logic fa_s5_c40_n13_s, fa_s5_c40_n13_c;
    logic fa_s5_c41_n14_s, fa_s5_c41_n14_c;
    logic fa_s5_c42_n15_s, fa_s5_c42_n15_c;
    logic fa_s5_c43_n16_s, fa_s5_c43_n16_c;
    logic fa_s5_c44_n17_s, fa_s5_c44_n17_c;
    logic fa_s5_c45_n18_s, fa_s5_c45_n18_c;
    logic fa_s5_c46_n19_s, fa_s5_c46_n19_c;
    logic fa_s5_c47_n20_s, fa_s5_c47_n20_c;
    logic fa_s5_c48_n21_s, fa_s5_c48_n21_c;
    logic fa_s5_c49_n22_s, fa_s5_c49_n22_c;
    logic fa_s5_c50_n23_s, fa_s5_c50_n23_c;
    logic fa_s5_c51_n24_s, fa_s5_c51_n24_c;
    logic fa_s5_c52_n25_s, fa_s5_c52_n25_c;
    logic fa_s5_c53_n26_s, fa_s5_c53_n26_c;
    logic fa_s5_c54_n27_s, fa_s5_c54_n27_c;
    logic fa_s5_c55_n28_s, fa_s5_c55_n28_c;
    logic fa_s5_c56_n29_s, fa_s5_c56_n29_c;
    logic fa_s5_c57_n30_s, fa_s5_c57_n30_c;
    logic fa_s5_c58_n31_s, fa_s5_c58_n31_c;
    logic fa_s5_c59_n32_s, fa_s5_c59_n32_c;
    logic fa_s5_c59_n33_s, fa_s5_c59_n33_c;
    logic fa_s5_c60_n34_s, fa_s5_c60_n34_c;
    logic fa_s5_c61_n35_s, fa_s5_c61_n35_c;
    logic fa_s5_c62_n36_s, fa_s5_c62_n36_c;
    logic fa_s5_c63_n37_s, fa_s5_c63_n37_c;
    logic fa_s5_c64_n38_s, fa_s5_c64_n38_c;
    logic fa_s5_c64_n39_s, fa_s5_c64_n39_c;
    logic fa_s5_c65_n40_s, fa_s5_c65_n40_c;
    logic fa_s5_c66_n41_s, fa_s5_c66_n41_c;
    logic fa_s5_c66_n42_s, fa_s5_c66_n42_c;
    logic fa_s5_c67_n43_s, fa_s5_c67_n43_c;
    logic fa_s5_c68_n44_s, fa_s5_c68_n44_c;
    logic fa_s5_c68_n45_s, fa_s5_c68_n45_c;
    logic fa_s5_c69_n46_s, fa_s5_c69_n46_c;
    logic fa_s5_c70_n47_s, fa_s5_c70_n47_c;
    logic fa_s5_c70_n48_s, fa_s5_c70_n48_c;
    logic fa_s5_c71_n49_s, fa_s5_c71_n49_c;
    logic fa_s5_c72_n50_s, fa_s5_c72_n50_c;
    logic fa_s5_c72_n51_s, fa_s5_c72_n51_c;
    logic fa_s5_c73_n52_s, fa_s5_c73_n52_c;
    logic fa_s5_c74_n53_s, fa_s5_c74_n53_c;
    logic fa_s5_c74_n54_s, fa_s5_c74_n54_c;
    logic fa_s5_c75_n55_s, fa_s5_c75_n55_c;
    logic fa_s5_c76_n56_s, fa_s5_c76_n56_c;
    logic fa_s5_c76_n57_s, fa_s5_c76_n57_c;
    logic fa_s5_c77_n58_s, fa_s5_c77_n58_c;
    logic fa_s5_c78_n59_s, fa_s5_c78_n59_c;
    logic fa_s5_c78_n60_s, fa_s5_c78_n60_c;
    logic fa_s5_c79_n61_s, fa_s5_c79_n61_c;
    logic fa_s5_c80_n62_s, fa_s5_c80_n62_c;
    logic fa_s5_c80_n63_s, fa_s5_c80_n63_c;
    logic fa_s5_c81_n64_s, fa_s5_c81_n64_c;
    logic fa_s5_c82_n65_s, fa_s5_c82_n65_c;
    logic fa_s5_c82_n66_s, fa_s5_c82_n66_c;
    logic fa_s5_c83_n67_s, fa_s5_c83_n67_c;
    logic fa_s5_c84_n68_s, fa_s5_c84_n68_c;
    logic fa_s5_c84_n69_s, fa_s5_c84_n69_c;
    logic fa_s5_c85_n70_s, fa_s5_c85_n70_c;
    logic fa_s5_c86_n71_s, fa_s5_c86_n71_c;
    logic fa_s5_c86_n72_s, fa_s5_c86_n72_c;
    logic fa_s5_c87_n73_s, fa_s5_c87_n73_c;
    logic fa_s5_c88_n74_s, fa_s5_c88_n74_c;
    logic fa_s5_c88_n75_s, fa_s5_c88_n75_c;
    logic fa_s5_c89_n76_s, fa_s5_c89_n76_c;
    logic fa_s5_c90_n77_s, fa_s5_c90_n77_c;
    logic fa_s5_c90_n78_s, fa_s5_c90_n78_c;
    logic fa_s5_c91_n79_s, fa_s5_c91_n79_c;
    logic fa_s5_c92_n80_s, fa_s5_c92_n80_c;
    logic fa_s5_c92_n81_s, fa_s5_c92_n81_c;
    logic fa_s5_c93_n82_s, fa_s5_c93_n82_c;
    logic fa_s5_c94_n83_s, fa_s5_c94_n83_c;
    logic fa_s5_c94_n84_s, fa_s5_c94_n84_c;
    logic fa_s5_c95_n85_s, fa_s5_c95_n85_c;
    logic fa_s5_c96_n86_s, fa_s5_c96_n86_c;
    logic fa_s5_c96_n87_s, fa_s5_c96_n87_c;
    logic fa_s5_c97_n88_s, fa_s5_c97_n88_c;
    logic fa_s5_c98_n89_s, fa_s5_c98_n89_c;
    logic fa_s5_c98_n90_s, fa_s5_c98_n90_c;
    logic fa_s5_c99_n91_s, fa_s5_c99_n91_c;
    logic fa_s5_c100_n92_s, fa_s5_c100_n92_c;
    logic fa_s5_c100_n93_s, fa_s5_c100_n93_c;
    logic fa_s5_c101_n94_s, fa_s5_c101_n94_c;
    logic fa_s5_c102_n95_s, fa_s5_c102_n95_c;
    logic fa_s5_c102_n96_s, fa_s5_c102_n96_c;
    logic fa_s5_c103_n97_s, fa_s5_c103_n97_c;
    logic fa_s5_c104_n98_s, fa_s5_c104_n98_c;
    logic fa_s5_c104_n99_s, fa_s5_c104_n99_c;
    logic fa_s5_c105_n100_s, fa_s5_c105_n100_c;
    logic fa_s5_c106_n101_s, fa_s5_c106_n101_c;
    logic fa_s5_c106_n102_s, fa_s5_c106_n102_c;
    logic fa_s5_c107_n103_s, fa_s5_c107_n103_c;
    logic fa_s5_c108_n104_s, fa_s5_c108_n104_c;
    logic fa_s5_c108_n105_s, fa_s5_c108_n105_c;
    logic fa_s5_c109_n106_s, fa_s5_c109_n106_c;
    logic fa_s5_c110_n107_s, fa_s5_c110_n107_c;
    logic fa_s5_c110_n108_s, fa_s5_c110_n108_c;
    logic fa_s5_c111_n109_s, fa_s5_c111_n109_c;
    logic fa_s5_c112_n110_s, fa_s5_c112_n110_c;
    logic fa_s5_c112_n111_s, fa_s5_c112_n111_c;
    logic fa_s5_c113_n112_s, fa_s5_c113_n112_c;
    logic fa_s5_c114_n113_s, fa_s5_c114_n113_c;
    logic fa_s5_c114_n114_s, fa_s5_c114_n114_c;
    logic fa_s5_c115_n115_s, fa_s5_c115_n115_c;
    logic fa_s5_c116_n116_s, fa_s5_c116_n116_c;
    logic fa_s5_c116_n117_s, fa_s5_c116_n117_c;
    logic fa_s5_c117_n118_s, fa_s5_c117_n118_c;
    logic fa_s5_c118_n119_s, fa_s5_c118_n119_c;
    logic fa_s5_c118_n120_s, fa_s5_c118_n120_c;
    logic fa_s5_c119_n121_s, fa_s5_c119_n121_c;
    logic fa_s5_c120_n122_s, fa_s5_c120_n122_c;
    logic fa_s5_c120_n123_s, fa_s5_c120_n123_c;
    logic fa_s5_c121_n124_s, fa_s5_c121_n124_c;
    logic fa_s5_c122_n125_s, fa_s5_c122_n125_c;
    logic fa_s5_c122_n126_s, fa_s5_c122_n126_c;
    logic fa_s5_c123_n127_s, fa_s5_c123_n127_c;
    logic fa_s5_c124_n128_s, fa_s5_c124_n128_c;
    logic fa_s5_c124_n129_s, fa_s5_c124_n129_c;
    logic fa_s5_c125_n130_s, fa_s5_c125_n130_c;
    logic fa_s5_c126_n131_s, fa_s5_c126_n131_c;
    logic fa_s5_c126_n132_s, fa_s5_c126_n132_c;
    logic fa_s6_c8_n0_s, fa_s6_c8_n0_c;
    logic fa_s6_c41_n1_s, fa_s6_c41_n1_c;
    logic fa_s6_c42_n2_s, fa_s6_c42_n2_c;
    logic fa_s6_c43_n3_s, fa_s6_c43_n3_c;
    logic fa_s6_c44_n4_s, fa_s6_c44_n4_c;
    logic fa_s6_c45_n5_s, fa_s6_c45_n5_c;
    logic fa_s6_c46_n6_s, fa_s6_c46_n6_c;
    logic fa_s6_c47_n7_s, fa_s6_c47_n7_c;
    logic fa_s6_c48_n8_s, fa_s6_c48_n8_c;
    logic fa_s6_c49_n9_s, fa_s6_c49_n9_c;
    logic fa_s6_c50_n10_s, fa_s6_c50_n10_c;
    logic fa_s6_c51_n11_s, fa_s6_c51_n11_c;
    logic fa_s6_c52_n12_s, fa_s6_c52_n12_c;
    logic fa_s6_c53_n13_s, fa_s6_c53_n13_c;
    logic fa_s6_c54_n14_s, fa_s6_c54_n14_c;
    logic fa_s6_c55_n15_s, fa_s6_c55_n15_c;
    logic fa_s6_c56_n16_s, fa_s6_c56_n16_c;
    logic fa_s6_c57_n17_s, fa_s6_c57_n17_c;
    logic fa_s6_c58_n18_s, fa_s6_c58_n18_c;
    logic fa_s6_c59_n19_s, fa_s6_c59_n19_c;
    logic fa_s6_c60_n20_s, fa_s6_c60_n20_c;
    logic fa_s6_c61_n21_s, fa_s6_c61_n21_c;
    logic fa_s6_c62_n22_s, fa_s6_c62_n22_c;
    logic fa_s6_c63_n23_s, fa_s6_c63_n23_c;
    logic fa_s6_c64_n24_s, fa_s6_c64_n24_c;
    logic fa_s6_c65_n25_s, fa_s6_c65_n25_c;
    logic fa_s6_c66_n26_s, fa_s6_c66_n26_c;
    logic fa_s6_c67_n27_s, fa_s6_c67_n27_c;
    logic fa_s6_c68_n28_s, fa_s6_c68_n28_c;
    logic fa_s6_c69_n29_s, fa_s6_c69_n29_c;
    logic fa_s6_c70_n30_s, fa_s6_c70_n30_c;
    logic fa_s6_c71_n31_s, fa_s6_c71_n31_c;
    logic fa_s6_c72_n32_s, fa_s6_c72_n32_c;
    logic fa_s6_c73_n33_s, fa_s6_c73_n33_c;
    logic fa_s6_c74_n34_s, fa_s6_c74_n34_c;
    logic fa_s6_c75_n35_s, fa_s6_c75_n35_c;
    logic fa_s6_c76_n36_s, fa_s6_c76_n36_c;
    logic fa_s6_c77_n37_s, fa_s6_c77_n37_c;
    logic fa_s6_c78_n38_s, fa_s6_c78_n38_c;
    logic fa_s6_c79_n39_s, fa_s6_c79_n39_c;
    logic fa_s6_c80_n40_s, fa_s6_c80_n40_c;
    logic fa_s6_c81_n41_s, fa_s6_c81_n41_c;
    logic fa_s6_c82_n42_s, fa_s6_c82_n42_c;
    logic fa_s6_c83_n43_s, fa_s6_c83_n43_c;
    logic fa_s6_c84_n44_s, fa_s6_c84_n44_c;
    logic fa_s6_c85_n45_s, fa_s6_c85_n45_c;
    logic fa_s6_c86_n46_s, fa_s6_c86_n46_c;
    logic fa_s6_c87_n47_s, fa_s6_c87_n47_c;
    logic fa_s6_c88_n48_s, fa_s6_c88_n48_c;
    logic fa_s6_c89_n49_s, fa_s6_c89_n49_c;
    logic fa_s6_c90_n50_s, fa_s6_c90_n50_c;
    logic fa_s6_c91_n51_s, fa_s6_c91_n51_c;
    logic fa_s6_c92_n52_s, fa_s6_c92_n52_c;
    logic fa_s6_c93_n53_s, fa_s6_c93_n53_c;
    logic fa_s6_c94_n54_s, fa_s6_c94_n54_c;
    logic fa_s6_c95_n55_s, fa_s6_c95_n55_c;
    logic fa_s6_c96_n56_s, fa_s6_c96_n56_c;
    logic fa_s6_c97_n57_s, fa_s6_c97_n57_c;
    logic fa_s6_c98_n58_s, fa_s6_c98_n58_c;
    logic fa_s6_c99_n59_s, fa_s6_c99_n59_c;
    logic fa_s6_c100_n60_s, fa_s6_c100_n60_c;
    logic fa_s6_c101_n61_s, fa_s6_c101_n61_c;
    logic fa_s6_c102_n62_s, fa_s6_c102_n62_c;
    logic fa_s6_c103_n63_s, fa_s6_c103_n63_c;
    logic fa_s6_c104_n64_s, fa_s6_c104_n64_c;
    logic fa_s6_c105_n65_s, fa_s6_c105_n65_c;
    logic fa_s6_c106_n66_s, fa_s6_c106_n66_c;
    logic fa_s6_c107_n67_s, fa_s6_c107_n67_c;
    logic fa_s6_c108_n68_s, fa_s6_c108_n68_c;
    logic fa_s6_c109_n69_s, fa_s6_c109_n69_c;
    logic fa_s6_c110_n70_s, fa_s6_c110_n70_c;
    logic fa_s6_c111_n71_s, fa_s6_c111_n71_c;
    logic fa_s6_c112_n72_s, fa_s6_c112_n72_c;
    logic fa_s6_c113_n73_s, fa_s6_c113_n73_c;
    logic fa_s6_c114_n74_s, fa_s6_c114_n74_c;
    logic fa_s6_c115_n75_s, fa_s6_c115_n75_c;
    logic fa_s6_c116_n76_s, fa_s6_c116_n76_c;
    logic fa_s6_c117_n77_s, fa_s6_c117_n77_c;
    logic fa_s6_c118_n78_s, fa_s6_c118_n78_c;
    logic fa_s6_c119_n79_s, fa_s6_c119_n79_c;
    logic fa_s6_c120_n80_s, fa_s6_c120_n80_c;
    logic fa_s6_c121_n81_s, fa_s6_c121_n81_c;
    logic fa_s6_c122_n82_s, fa_s6_c122_n82_c;
    logic fa_s6_c123_n83_s, fa_s6_c123_n83_c;
    logic fa_s6_c124_n84_s, fa_s6_c124_n84_c;
    logic fa_s6_c125_n85_s, fa_s6_c125_n85_c;
    logic fa_s6_c126_n86_s, fa_s6_c126_n86_c;
    logic fa_s7_c9_n0_s, fa_s7_c9_n0_c;
    logic fa_s7_c60_n1_s, fa_s7_c60_n1_c;
    logic fa_s7_c61_n2_s, fa_s7_c61_n2_c;
    logic fa_s7_c62_n3_s, fa_s7_c62_n3_c;
    logic fa_s7_c63_n4_s, fa_s7_c63_n4_c;
    logic fa_s7_c64_n5_s, fa_s7_c64_n5_c;
    logic fa_s7_c65_n6_s, fa_s7_c65_n6_c;
    logic fa_s7_c66_n7_s, fa_s7_c66_n7_c;
    logic fa_s7_c67_n8_s, fa_s7_c67_n8_c;
    logic fa_s7_c68_n9_s, fa_s7_c68_n9_c;
    logic fa_s7_c69_n10_s, fa_s7_c69_n10_c;
    logic fa_s7_c70_n11_s, fa_s7_c70_n11_c;
    logic fa_s7_c71_n12_s, fa_s7_c71_n12_c;
    logic fa_s7_c72_n13_s, fa_s7_c72_n13_c;
    logic fa_s7_c73_n14_s, fa_s7_c73_n14_c;
    logic fa_s7_c74_n15_s, fa_s7_c74_n15_c;
    logic fa_s7_c75_n16_s, fa_s7_c75_n16_c;
    logic fa_s7_c76_n17_s, fa_s7_c76_n17_c;
    logic fa_s7_c77_n18_s, fa_s7_c77_n18_c;
    logic fa_s7_c78_n19_s, fa_s7_c78_n19_c;
    logic fa_s7_c79_n20_s, fa_s7_c79_n20_c;
    logic fa_s7_c80_n21_s, fa_s7_c80_n21_c;
    logic fa_s7_c81_n22_s, fa_s7_c81_n22_c;
    logic fa_s7_c82_n23_s, fa_s7_c82_n23_c;
    logic fa_s7_c83_n24_s, fa_s7_c83_n24_c;
    logic fa_s7_c84_n25_s, fa_s7_c84_n25_c;
    logic fa_s7_c85_n26_s, fa_s7_c85_n26_c;
    logic fa_s7_c86_n27_s, fa_s7_c86_n27_c;
    logic fa_s7_c87_n28_s, fa_s7_c87_n28_c;
    logic fa_s7_c88_n29_s, fa_s7_c88_n29_c;
    logic fa_s7_c89_n30_s, fa_s7_c89_n30_c;
    logic fa_s7_c90_n31_s, fa_s7_c90_n31_c;
    logic fa_s7_c91_n32_s, fa_s7_c91_n32_c;
    logic fa_s7_c92_n33_s, fa_s7_c92_n33_c;
    logic fa_s7_c93_n34_s, fa_s7_c93_n34_c;
    logic fa_s7_c94_n35_s, fa_s7_c94_n35_c;
    logic fa_s7_c95_n36_s, fa_s7_c95_n36_c;
    logic fa_s7_c96_n37_s, fa_s7_c96_n37_c;
    logic fa_s7_c97_n38_s, fa_s7_c97_n38_c;
    logic fa_s7_c98_n39_s, fa_s7_c98_n39_c;
    logic fa_s7_c99_n40_s, fa_s7_c99_n40_c;
    logic fa_s7_c100_n41_s, fa_s7_c100_n41_c;
    logic fa_s7_c101_n42_s, fa_s7_c101_n42_c;
    logic fa_s7_c102_n43_s, fa_s7_c102_n43_c;
    logic fa_s7_c103_n44_s, fa_s7_c103_n44_c;
    logic fa_s7_c104_n45_s, fa_s7_c104_n45_c;
    logic fa_s7_c105_n46_s, fa_s7_c105_n46_c;
    logic fa_s7_c106_n47_s, fa_s7_c106_n47_c;
    logic fa_s7_c107_n48_s, fa_s7_c107_n48_c;
    logic fa_s7_c108_n49_s, fa_s7_c108_n49_c;
    logic fa_s7_c109_n50_s, fa_s7_c109_n50_c;
    logic fa_s7_c110_n51_s, fa_s7_c110_n51_c;
    logic fa_s7_c111_n52_s, fa_s7_c111_n52_c;
    logic fa_s7_c112_n53_s, fa_s7_c112_n53_c;
    logic fa_s7_c113_n54_s, fa_s7_c113_n54_c;
    logic fa_s7_c114_n55_s, fa_s7_c114_n55_c;
    logic fa_s7_c115_n56_s, fa_s7_c115_n56_c;
    logic fa_s7_c116_n57_s, fa_s7_c116_n57_c;
    logic fa_s7_c117_n58_s, fa_s7_c117_n58_c;
    logic fa_s7_c118_n59_s, fa_s7_c118_n59_c;
    logic fa_s7_c119_n60_s, fa_s7_c119_n60_c;
    logic fa_s7_c120_n61_s, fa_s7_c120_n61_c;
    logic fa_s7_c121_n62_s, fa_s7_c121_n62_c;
    logic fa_s7_c122_n63_s, fa_s7_c122_n63_c;
    logic fa_s7_c123_n64_s, fa_s7_c123_n64_c;
    logic fa_s7_c124_n65_s, fa_s7_c124_n65_c;
    logic fa_s7_c125_n66_s, fa_s7_c125_n66_c;
    logic fa_s7_c126_n67_s, fa_s7_c126_n67_c;
    logic ha_s0_c0_n0_s, ha_s0_c0_n0_c;
    logic ha_s1_c1_n0_s, ha_s1_c1_n0_c;
    logic ha_s2_c2_n0_s, ha_s2_c2_n0_c;
    logic ha_s3_c3_n0_s, ha_s3_c3_n0_c;
    logic ha_s4_c4_n0_s, ha_s4_c4_n0_c;
    logic ha_s5_c5_n0_s, ha_s5_c5_n0_c;
    logic ha_s5_c60_n1_s, ha_s5_c60_n1_c;
    logic ha_s5_c61_n2_s, ha_s5_c61_n2_c;
    logic ha_s5_c62_n3_s, ha_s5_c62_n3_c;
    logic ha_s5_c63_n4_s, ha_s5_c63_n4_c;
    logic ha_s5_c65_n5_s, ha_s5_c65_n5_c;
    logic ha_s5_c67_n6_s, ha_s5_c67_n6_c;
    logic ha_s5_c69_n7_s, ha_s5_c69_n7_c;
    logic ha_s5_c71_n8_s, ha_s5_c71_n8_c;
    logic ha_s5_c73_n9_s, ha_s5_c73_n9_c;
    logic ha_s5_c75_n10_s, ha_s5_c75_n10_c;
    logic ha_s5_c77_n11_s, ha_s5_c77_n11_c;
    logic ha_s5_c79_n12_s, ha_s5_c79_n12_c;
    logic ha_s5_c81_n13_s, ha_s5_c81_n13_c;
    logic ha_s5_c83_n14_s, ha_s5_c83_n14_c;
    logic ha_s5_c85_n15_s, ha_s5_c85_n15_c;
    logic ha_s5_c87_n16_s, ha_s5_c87_n16_c;
    logic ha_s5_c89_n17_s, ha_s5_c89_n17_c;
    logic ha_s5_c91_n18_s, ha_s5_c91_n18_c;
    logic ha_s5_c93_n19_s, ha_s5_c93_n19_c;
    logic ha_s5_c95_n20_s, ha_s5_c95_n20_c;
    logic ha_s5_c97_n21_s, ha_s5_c97_n21_c;
    logic ha_s5_c99_n22_s, ha_s5_c99_n22_c;
    logic ha_s5_c101_n23_s, ha_s5_c101_n23_c;
    logic ha_s5_c103_n24_s, ha_s5_c103_n24_c;
    logic ha_s5_c105_n25_s, ha_s5_c105_n25_c;
    logic ha_s5_c107_n26_s, ha_s5_c107_n26_c;
    logic ha_s5_c109_n27_s, ha_s5_c109_n27_c;
    logic ha_s5_c111_n28_s, ha_s5_c111_n28_c;
    logic ha_s5_c113_n29_s, ha_s5_c113_n29_c;
    logic ha_s5_c115_n30_s, ha_s5_c115_n30_c;
    logic ha_s5_c117_n31_s, ha_s5_c117_n31_c;
    logic ha_s5_c119_n32_s, ha_s5_c119_n32_c;
    logic ha_s5_c121_n33_s, ha_s5_c121_n33_c;
    logic ha_s5_c123_n34_s, ha_s5_c123_n34_c;
    logic ha_s5_c125_n35_s, ha_s5_c125_n35_c;
    logic ha_s6_c6_n0_s, ha_s6_c6_n0_c;
    logic ha_s7_c7_n0_s, ha_s7_c7_n0_c;
    logic ha_s7_c10_n1_s, ha_s7_c10_n1_c;
    logic ha_s7_c11_n2_s, ha_s7_c11_n2_c;
    logic ha_s7_c12_n3_s, ha_s7_c12_n3_c;
    logic ha_s7_c13_n4_s, ha_s7_c13_n4_c;
    logic ha_s7_c14_n5_s, ha_s7_c14_n5_c;
    logic ha_s7_c15_n6_s, ha_s7_c15_n6_c;
    logic ha_s7_c16_n7_s, ha_s7_c16_n7_c;
    logic ha_s7_c17_n8_s, ha_s7_c17_n8_c;
    logic ha_s7_c18_n9_s, ha_s7_c18_n9_c;
    logic ha_s7_c19_n10_s, ha_s7_c19_n10_c;
    logic ha_s7_c20_n11_s, ha_s7_c20_n11_c;
    logic ha_s7_c21_n12_s, ha_s7_c21_n12_c;
    logic ha_s7_c22_n13_s, ha_s7_c22_n13_c;
    logic ha_s7_c23_n14_s, ha_s7_c23_n14_c;
    logic ha_s7_c24_n15_s, ha_s7_c24_n15_c;
    logic ha_s7_c25_n16_s, ha_s7_c25_n16_c;
    logic ha_s7_c26_n17_s, ha_s7_c26_n17_c;
    logic ha_s7_c27_n18_s, ha_s7_c27_n18_c;
    logic ha_s7_c28_n19_s, ha_s7_c28_n19_c;
    logic ha_s7_c29_n20_s, ha_s7_c29_n20_c;
    logic ha_s7_c30_n21_s, ha_s7_c30_n21_c;
    logic ha_s7_c31_n22_s, ha_s7_c31_n22_c;
    logic ha_s7_c32_n23_s, ha_s7_c32_n23_c;
    logic ha_s7_c33_n24_s, ha_s7_c33_n24_c;
    logic ha_s7_c34_n25_s, ha_s7_c34_n25_c;
    logic ha_s7_c35_n26_s, ha_s7_c35_n26_c;
    logic ha_s7_c36_n27_s, ha_s7_c36_n27_c;
    logic ha_s7_c37_n28_s, ha_s7_c37_n28_c;
    logic ha_s7_c38_n29_s, ha_s7_c38_n29_c;
    logic ha_s7_c39_n30_s, ha_s7_c39_n30_c;
    logic ha_s7_c40_n31_s, ha_s7_c40_n31_c;
    logic ha_s7_c41_n32_s, ha_s7_c41_n32_c;
    logic ha_s7_c42_n33_s, ha_s7_c42_n33_c;
    logic ha_s7_c43_n34_s, ha_s7_c43_n34_c;
    logic ha_s7_c44_n35_s, ha_s7_c44_n35_c;
    logic ha_s7_c45_n36_s, ha_s7_c45_n36_c;
    logic ha_s7_c46_n37_s, ha_s7_c46_n37_c;
    logic ha_s7_c47_n38_s, ha_s7_c47_n38_c;
    logic ha_s7_c48_n39_s, ha_s7_c48_n39_c;
    logic ha_s7_c49_n40_s, ha_s7_c49_n40_c;
    logic ha_s7_c50_n41_s, ha_s7_c50_n41_c;
    logic ha_s7_c51_n42_s, ha_s7_c51_n42_c;
    logic ha_s7_c52_n43_s, ha_s7_c52_n43_c;
    logic ha_s7_c53_n44_s, ha_s7_c53_n44_c;
    logic ha_s7_c54_n45_s, ha_s7_c54_n45_c;
    logic ha_s7_c55_n46_s, ha_s7_c55_n46_c;
    logic ha_s7_c56_n47_s, ha_s7_c56_n47_c;
    logic ha_s7_c57_n48_s, ha_s7_c57_n48_c;
    logic ha_s7_c58_n49_s, ha_s7_c58_n49_c;
    logic ha_s7_c59_n50_s, ha_s7_c59_n50_c;

    // Stage 0 signals
    logic [1:0] stage0_col0;
    logic [0:0] stage0_col1;
    logic [2:0] stage0_col2;
    logic [1:0] stage0_col3;
    logic [3:0] stage0_col4;
    logic [2:0] stage0_col5;
    logic [4:0] stage0_col6;
    logic [3:0] stage0_col7;
    logic [5:0] stage0_col8;
    logic [4:0] stage0_col9;
    logic [6:0] stage0_col10;
    logic [5:0] stage0_col11;
    logic [7:0] stage0_col12;
    logic [6:0] stage0_col13;
    logic [8:0] stage0_col14;
    logic [7:0] stage0_col15;
    logic [9:0] stage0_col16;
    logic [8:0] stage0_col17;
    logic [10:0] stage0_col18;
    logic [9:0] stage0_col19;
    logic [11:0] stage0_col20;
    logic [10:0] stage0_col21;
    logic [12:0] stage0_col22;
    logic [11:0] stage0_col23;
    logic [13:0] stage0_col24;
    logic [12:0] stage0_col25;
    logic [14:0] stage0_col26;
    logic [13:0] stage0_col27;
    logic [15:0] stage0_col28;
    logic [14:0] stage0_col29;
    logic [16:0] stage0_col30;
    logic [15:0] stage0_col31;
    logic [17:0] stage0_col32;
    logic [16:0] stage0_col33;
    logic [18:0] stage0_col34;
    logic [17:0] stage0_col35;
    logic [19:0] stage0_col36;
    logic [18:0] stage0_col37;
    logic [20:0] stage0_col38;
    logic [19:0] stage0_col39;
    logic [21:0] stage0_col40;
    logic [20:0] stage0_col41;
    logic [22:0] stage0_col42;
    logic [21:0] stage0_col43;
    logic [23:0] stage0_col44;
    logic [22:0] stage0_col45;
    logic [24:0] stage0_col46;
    logic [23:0] stage0_col47;
    logic [25:0] stage0_col48;
    logic [24:0] stage0_col49;
    logic [26:0] stage0_col50;
    logic [25:0] stage0_col51;
    logic [27:0] stage0_col52;
    logic [26:0] stage0_col53;
    logic [28:0] stage0_col54;
    logic [27:0] stage0_col55;
    logic [29:0] stage0_col56;
    logic [28:0] stage0_col57;
    logic [30:0] stage0_col58;
    logic [29:0] stage0_col59;
    logic [31:0] stage0_col60;
    logic [30:0] stage0_col61;
    logic [32:0] stage0_col62;
    logic [31:0] stage0_col63;
    logic [32:0] stage0_col64;
    logic [31:0] stage0_col65;
    logic [32:0] stage0_col66;
    logic [31:0] stage0_col67;
    logic [32:0] stage0_col68;
    logic [31:0] stage0_col69;
    logic [32:0] stage0_col70;
    logic [31:0] stage0_col71;
    logic [32:0] stage0_col72;
    logic [31:0] stage0_col73;
    logic [32:0] stage0_col74;
    logic [31:0] stage0_col75;
    logic [32:0] stage0_col76;
    logic [31:0] stage0_col77;
    logic [32:0] stage0_col78;
    logic [31:0] stage0_col79;
    logic [32:0] stage0_col80;
    logic [31:0] stage0_col81;
    logic [32:0] stage0_col82;
    logic [31:0] stage0_col83;
    logic [32:0] stage0_col84;
    logic [31:0] stage0_col85;
    logic [32:0] stage0_col86;
    logic [31:0] stage0_col87;
    logic [32:0] stage0_col88;
    logic [31:0] stage0_col89;
    logic [32:0] stage0_col90;
    logic [31:0] stage0_col91;
    logic [32:0] stage0_col92;
    logic [31:0] stage0_col93;
    logic [32:0] stage0_col94;
    logic [31:0] stage0_col95;
    logic [32:0] stage0_col96;
    logic [31:0] stage0_col97;
    logic [32:0] stage0_col98;
    logic [31:0] stage0_col99;
    logic [32:0] stage0_col100;
    logic [31:0] stage0_col101;
    logic [32:0] stage0_col102;
    logic [31:0] stage0_col103;
    logic [32:0] stage0_col104;
    logic [31:0] stage0_col105;
    logic [32:0] stage0_col106;
    logic [31:0] stage0_col107;
    logic [32:0] stage0_col108;
    logic [31:0] stage0_col109;
    logic [32:0] stage0_col110;
    logic [31:0] stage0_col111;
    logic [32:0] stage0_col112;
    logic [31:0] stage0_col113;
    logic [32:0] stage0_col114;
    logic [31:0] stage0_col115;
    logic [32:0] stage0_col116;
    logic [31:0] stage0_col117;
    logic [32:0] stage0_col118;
    logic [31:0] stage0_col119;
    logic [32:0] stage0_col120;
    logic [31:0] stage0_col121;
    logic [32:0] stage0_col122;
    logic [31:0] stage0_col123;
    logic [32:0] stage0_col124;
    logic [31:0] stage0_col125;
    logic [32:0] stage0_col126;
    logic [31:0] stage0_col127;

    // Stage 1 signals
    logic [0:0] stage1_col0;
    logic [1:0] stage1_col1;
    logic [0:0] stage1_col2;
    logic [2:0] stage1_col3;
    logic [1:0] stage1_col4;
    logic [1:0] stage1_col5;
    logic [3:0] stage1_col6;
    logic [2:0] stage1_col7;
    logic [2:0] stage1_col8;
    logic [4:0] stage1_col9;
    logic [3:0] stage1_col10;
    logic [3:0] stage1_col11;
    logic [5:0] stage1_col12;
    logic [4:0] stage1_col13;
    logic [4:0] stage1_col14;
    logic [6:0] stage1_col15;
    logic [5:0] stage1_col16;
    logic [5:0] stage1_col17;
    logic [7:0] stage1_col18;
    logic [6:0] stage1_col19;
    logic [6:0] stage1_col20;
    logic [8:0] stage1_col21;
    logic [7:0] stage1_col22;
    logic [7:0] stage1_col23;
    logic [9:0] stage1_col24;
    logic [8:0] stage1_col25;
    logic [8:0] stage1_col26;
    logic [10:0] stage1_col27;
    logic [9:0] stage1_col28;
    logic [9:0] stage1_col29;
    logic [11:0] stage1_col30;
    logic [10:0] stage1_col31;
    logic [10:0] stage1_col32;
    logic [12:0] stage1_col33;
    logic [11:0] stage1_col34;
    logic [11:0] stage1_col35;
    logic [13:0] stage1_col36;
    logic [12:0] stage1_col37;
    logic [12:0] stage1_col38;
    logic [14:0] stage1_col39;
    logic [13:0] stage1_col40;
    logic [13:0] stage1_col41;
    logic [15:0] stage1_col42;
    logic [14:0] stage1_col43;
    logic [14:0] stage1_col44;
    logic [16:0] stage1_col45;
    logic [15:0] stage1_col46;
    logic [15:0] stage1_col47;
    logic [17:0] stage1_col48;
    logic [16:0] stage1_col49;
    logic [16:0] stage1_col50;
    logic [18:0] stage1_col51;
    logic [17:0] stage1_col52;
    logic [17:0] stage1_col53;
    logic [19:0] stage1_col54;
    logic [18:0] stage1_col55;
    logic [18:0] stage1_col56;
    logic [20:0] stage1_col57;
    logic [19:0] stage1_col58;
    logic [19:0] stage1_col59;
    logic [21:0] stage1_col60;
    logic [20:0] stage1_col61;
    logic [20:0] stage1_col62;
    logic [22:0] stage1_col63;
    logic [20:0] stage1_col64;
    logic [22:0] stage1_col65;
    logic [20:0] stage1_col66;
    logic [22:0] stage1_col67;
    logic [20:0] stage1_col68;
    logic [22:0] stage1_col69;
    logic [20:0] stage1_col70;
    logic [22:0] stage1_col71;
    logic [20:0] stage1_col72;
    logic [22:0] stage1_col73;
    logic [20:0] stage1_col74;
    logic [22:0] stage1_col75;
    logic [20:0] stage1_col76;
    logic [22:0] stage1_col77;
    logic [20:0] stage1_col78;
    logic [22:0] stage1_col79;
    logic [20:0] stage1_col80;
    logic [22:0] stage1_col81;
    logic [20:0] stage1_col82;
    logic [22:0] stage1_col83;
    logic [20:0] stage1_col84;
    logic [22:0] stage1_col85;
    logic [20:0] stage1_col86;
    logic [22:0] stage1_col87;
    logic [20:0] stage1_col88;
    logic [22:0] stage1_col89;
    logic [20:0] stage1_col90;
    logic [22:0] stage1_col91;
    logic [20:0] stage1_col92;
    logic [22:0] stage1_col93;
    logic [20:0] stage1_col94;
    logic [22:0] stage1_col95;
    logic [20:0] stage1_col96;
    logic [22:0] stage1_col97;
    logic [20:0] stage1_col98;
    logic [22:0] stage1_col99;
    logic [20:0] stage1_col100;
    logic [22:0] stage1_col101;
    logic [20:0] stage1_col102;
    logic [22:0] stage1_col103;
    logic [20:0] stage1_col104;
    logic [22:0] stage1_col105;
    logic [20:0] stage1_col106;
    logic [22:0] stage1_col107;
    logic [20:0] stage1_col108;
    logic [22:0] stage1_col109;
    logic [20:0] stage1_col110;
    logic [22:0] stage1_col111;
    logic [20:0] stage1_col112;
    logic [22:0] stage1_col113;
    logic [20:0] stage1_col114;
    logic [22:0] stage1_col115;
    logic [20:0] stage1_col116;
    logic [22:0] stage1_col117;
    logic [20:0] stage1_col118;
    logic [22:0] stage1_col119;
    logic [20:0] stage1_col120;
    logic [22:0] stage1_col121;
    logic [20:0] stage1_col122;
    logic [22:0] stage1_col123;
    logic [20:0] stage1_col124;
    logic [22:0] stage1_col125;
    logic [20:0] stage1_col126;
    logic [42:0] stage1_col127;

    // Stage 2 signals
    logic [0:0] stage2_col0;
    logic [0:0] stage2_col1;
    logic [1:0] stage2_col2;
    logic [0:0] stage2_col3;
    logic [2:0] stage2_col4;
    logic [1:0] stage2_col5;
    logic [1:0] stage2_col6;
    logic [1:0] stage2_col7;
    logic [1:0] stage2_col8;
    logic [3:0] stage2_col9;
    logic [2:0] stage2_col10;
    logic [2:0] stage2_col11;
    logic [2:0] stage2_col12;
    logic [4:0] stage2_col13;
    logic [3:0] stage2_col14;
    logic [3:0] stage2_col15;
    logic [3:0] stage2_col16;
    logic [3:0] stage2_col17;
    logic [5:0] stage2_col18;
    logic [4:0] stage2_col19;
    logic [4:0] stage2_col20;
    logic [4:0] stage2_col21;
    logic [6:0] stage2_col22;
    logic [5:0] stage2_col23;
    logic [5:0] stage2_col24;
    logic [5:0] stage2_col25;
    logic [5:0] stage2_col26;
    logic [7:0] stage2_col27;
    logic [6:0] stage2_col28;
    logic [6:0] stage2_col29;
    logic [6:0] stage2_col30;
    logic [8:0] stage2_col31;
    logic [7:0] stage2_col32;
    logic [7:0] stage2_col33;
    logic [7:0] stage2_col34;
    logic [7:0] stage2_col35;
    logic [9:0] stage2_col36;
    logic [8:0] stage2_col37;
    logic [8:0] stage2_col38;
    logic [8:0] stage2_col39;
    logic [10:0] stage2_col40;
    logic [9:0] stage2_col41;
    logic [9:0] stage2_col42;
    logic [9:0] stage2_col43;
    logic [9:0] stage2_col44;
    logic [11:0] stage2_col45;
    logic [10:0] stage2_col46;
    logic [10:0] stage2_col47;
    logic [10:0] stage2_col48;
    logic [12:0] stage2_col49;
    logic [11:0] stage2_col50;
    logic [11:0] stage2_col51;
    logic [11:0] stage2_col52;
    logic [11:0] stage2_col53;
    logic [13:0] stage2_col54;
    logic [12:0] stage2_col55;
    logic [12:0] stage2_col56;
    logic [12:0] stage2_col57;
    logic [14:0] stage2_col58;
    logic [13:0] stage2_col59;
    logic [13:0] stage2_col60;
    logic [13:0] stage2_col61;
    logic [13:0] stage2_col62;
    logic [15:0] stage2_col63;
    logic [13:0] stage2_col64;
    logic [15:0] stage2_col65;
    logic [13:0] stage2_col66;
    logic [15:0] stage2_col67;
    logic [13:0] stage2_col68;
    logic [15:0] stage2_col69;
    logic [13:0] stage2_col70;
    logic [15:0] stage2_col71;
    logic [13:0] stage2_col72;
    logic [15:0] stage2_col73;
    logic [13:0] stage2_col74;
    logic [15:0] stage2_col75;
    logic [13:0] stage2_col76;
    logic [15:0] stage2_col77;
    logic [13:0] stage2_col78;
    logic [15:0] stage2_col79;
    logic [13:0] stage2_col80;
    logic [15:0] stage2_col81;
    logic [13:0] stage2_col82;
    logic [15:0] stage2_col83;
    logic [13:0] stage2_col84;
    logic [15:0] stage2_col85;
    logic [13:0] stage2_col86;
    logic [15:0] stage2_col87;
    logic [13:0] stage2_col88;
    logic [15:0] stage2_col89;
    logic [13:0] stage2_col90;
    logic [15:0] stage2_col91;
    logic [13:0] stage2_col92;
    logic [15:0] stage2_col93;
    logic [13:0] stage2_col94;
    logic [15:0] stage2_col95;
    logic [13:0] stage2_col96;
    logic [15:0] stage2_col97;
    logic [13:0] stage2_col98;
    logic [15:0] stage2_col99;
    logic [13:0] stage2_col100;
    logic [15:0] stage2_col101;
    logic [13:0] stage2_col102;
    logic [15:0] stage2_col103;
    logic [13:0] stage2_col104;
    logic [15:0] stage2_col105;
    logic [13:0] stage2_col106;
    logic [15:0] stage2_col107;
    logic [13:0] stage2_col108;
    logic [15:0] stage2_col109;
    logic [13:0] stage2_col110;
    logic [15:0] stage2_col111;
    logic [13:0] stage2_col112;
    logic [15:0] stage2_col113;
    logic [13:0] stage2_col114;
    logic [15:0] stage2_col115;
    logic [13:0] stage2_col116;
    logic [15:0] stage2_col117;
    logic [13:0] stage2_col118;
    logic [15:0] stage2_col119;
    logic [13:0] stage2_col120;
    logic [15:0] stage2_col121;
    logic [13:0] stage2_col122;
    logic [15:0] stage2_col123;
    logic [13:0] stage2_col124;
    logic [15:0] stage2_col125;
    logic [13:0] stage2_col126;
    logic [49:0] stage2_col127;

    // Stage 3 signals
    logic [0:0] stage3_col0;
    logic [0:0] stage3_col1;
    logic [0:0] stage3_col2;
    logic [1:0] stage3_col3;
    logic [0:0] stage3_col4;
    logic [2:0] stage3_col5;
    logic [1:0] stage3_col6;
    logic [1:0] stage3_col7;
    logic [1:0] stage3_col8;
    logic [1:0] stage3_col9;
    logic [1:0] stage3_col10;
    logic [1:0] stage3_col11;
    logic [1:0] stage3_col12;
    logic [3:0] stage3_col13;
    logic [2:0] stage3_col14;
    logic [2:0] stage3_col15;
    logic [2:0] stage3_col16;
    logic [2:0] stage3_col17;
    logic [2:0] stage3_col18;
    logic [4:0] stage3_col19;
    logic [3:0] stage3_col20;
    logic [3:0] stage3_col21;
    logic [3:0] stage3_col22;
    logic [3:0] stage3_col23;
    logic [3:0] stage3_col24;
    logic [3:0] stage3_col25;
    logic [3:0] stage3_col26;
    logic [5:0] stage3_col27;
    logic [4:0] stage3_col28;
    logic [4:0] stage3_col29;
    logic [4:0] stage3_col30;
    logic [4:0] stage3_col31;
    logic [6:0] stage3_col32;
    logic [5:0] stage3_col33;
    logic [5:0] stage3_col34;
    logic [5:0] stage3_col35;
    logic [5:0] stage3_col36;
    logic [5:0] stage3_col37;
    logic [5:0] stage3_col38;
    logic [5:0] stage3_col39;
    logic [7:0] stage3_col40;
    logic [6:0] stage3_col41;
    logic [6:0] stage3_col42;
    logic [6:0] stage3_col43;
    logic [6:0] stage3_col44;
    logic [6:0] stage3_col45;
    logic [8:0] stage3_col46;
    logic [7:0] stage3_col47;
    logic [7:0] stage3_col48;
    logic [7:0] stage3_col49;
    logic [7:0] stage3_col50;
    logic [7:0] stage3_col51;
    logic [7:0] stage3_col52;
    logic [7:0] stage3_col53;
    logic [9:0] stage3_col54;
    logic [8:0] stage3_col55;
    logic [8:0] stage3_col56;
    logic [8:0] stage3_col57;
    logic [8:0] stage3_col58;
    logic [10:0] stage3_col59;
    logic [9:0] stage3_col60;
    logic [9:0] stage3_col61;
    logic [9:0] stage3_col62;
    logic [9:0] stage3_col63;
    logic [10:0] stage3_col64;
    logic [9:0] stage3_col65;
    logic [10:0] stage3_col66;
    logic [9:0] stage3_col67;
    logic [10:0] stage3_col68;
    logic [9:0] stage3_col69;
    logic [10:0] stage3_col70;
    logic [9:0] stage3_col71;
    logic [10:0] stage3_col72;
    logic [9:0] stage3_col73;
    logic [10:0] stage3_col74;
    logic [9:0] stage3_col75;
    logic [10:0] stage3_col76;
    logic [9:0] stage3_col77;
    logic [10:0] stage3_col78;
    logic [9:0] stage3_col79;
    logic [10:0] stage3_col80;
    logic [9:0] stage3_col81;
    logic [10:0] stage3_col82;
    logic [9:0] stage3_col83;
    logic [10:0] stage3_col84;
    logic [9:0] stage3_col85;
    logic [10:0] stage3_col86;
    logic [9:0] stage3_col87;
    logic [10:0] stage3_col88;
    logic [9:0] stage3_col89;
    logic [10:0] stage3_col90;
    logic [9:0] stage3_col91;
    logic [10:0] stage3_col92;
    logic [9:0] stage3_col93;
    logic [10:0] stage3_col94;
    logic [9:0] stage3_col95;
    logic [10:0] stage3_col96;
    logic [9:0] stage3_col97;
    logic [10:0] stage3_col98;
    logic [9:0] stage3_col99;
    logic [10:0] stage3_col100;
    logic [9:0] stage3_col101;
    logic [10:0] stage3_col102;
    logic [9:0] stage3_col103;
    logic [10:0] stage3_col104;
    logic [9:0] stage3_col105;
    logic [10:0] stage3_col106;
    logic [9:0] stage3_col107;
    logic [10:0] stage3_col108;
    logic [9:0] stage3_col109;
    logic [10:0] stage3_col110;
    logic [9:0] stage3_col111;
    logic [10:0] stage3_col112;
    logic [9:0] stage3_col113;
    logic [10:0] stage3_col114;
    logic [9:0] stage3_col115;
    logic [10:0] stage3_col116;
    logic [9:0] stage3_col117;
    logic [10:0] stage3_col118;
    logic [9:0] stage3_col119;
    logic [10:0] stage3_col120;
    logic [9:0] stage3_col121;
    logic [10:0] stage3_col122;
    logic [9:0] stage3_col123;
    logic [10:0] stage3_col124;
    logic [9:0] stage3_col125;
    logic [10:0] stage3_col126;
    logic [53:0] stage3_col127;

    // Stage 4 signals
    logic [0:0] stage4_col0;
    logic [0:0] stage4_col1;
    logic [0:0] stage4_col2;
    logic [0:0] stage4_col3;
    logic [1:0] stage4_col4;
    logic [0:0] stage4_col5;
    logic [2:0] stage4_col6;
    logic [1:0] stage4_col7;
    logic [1:0] stage4_col8;
    logic [1:0] stage4_col9;
    logic [1:0] stage4_col10;
    logic [1:0] stage4_col11;
    logic [1:0] stage4_col12;
    logic [1:0] stage4_col13;
    logic [1:0] stage4_col14;
    logic [1:0] stage4_col15;
    logic [1:0] stage4_col16;
    logic [1:0] stage4_col17;
    logic [1:0] stage4_col18;
    logic [3:0] stage4_col19;
    logic [2:0] stage4_col20;
    logic [2:0] stage4_col21;
    logic [2:0] stage4_col22;
    logic [2:0] stage4_col23;
    logic [2:0] stage4_col24;
    logic [2:0] stage4_col25;
    logic [2:0] stage4_col26;
    logic [2:0] stage4_col27;
    logic [4:0] stage4_col28;
    logic [3:0] stage4_col29;
    logic [3:0] stage4_col30;
    logic [3:0] stage4_col31;
    logic [3:0] stage4_col32;
    logic [3:0] stage4_col33;
    logic [3:0] stage4_col34;
    logic [3:0] stage4_col35;
    logic [3:0] stage4_col36;
    logic [3:0] stage4_col37;
    logic [3:0] stage4_col38;
    logic [3:0] stage4_col39;
    logic [5:0] stage4_col40;
    logic [4:0] stage4_col41;
    logic [4:0] stage4_col42;
    logic [4:0] stage4_col43;
    logic [4:0] stage4_col44;
    logic [4:0] stage4_col45;
    logic [4:0] stage4_col46;
    logic [6:0] stage4_col47;
    logic [5:0] stage4_col48;
    logic [5:0] stage4_col49;
    logic [5:0] stage4_col50;
    logic [5:0] stage4_col51;
    logic [5:0] stage4_col52;
    logic [5:0] stage4_col53;
    logic [5:0] stage4_col54;
    logic [5:0] stage4_col55;
    logic [5:0] stage4_col56;
    logic [5:0] stage4_col57;
    logic [5:0] stage4_col58;
    logic [7:0] stage4_col59;
    logic [6:0] stage4_col60;
    logic [6:0] stage4_col61;
    logic [6:0] stage4_col62;
    logic [6:0] stage4_col63;
    logic [7:0] stage4_col64;
    logic [6:0] stage4_col65;
    logic [7:0] stage4_col66;
    logic [6:0] stage4_col67;
    logic [7:0] stage4_col68;
    logic [6:0] stage4_col69;
    logic [7:0] stage4_col70;
    logic [6:0] stage4_col71;
    logic [7:0] stage4_col72;
    logic [6:0] stage4_col73;
    logic [7:0] stage4_col74;
    logic [6:0] stage4_col75;
    logic [7:0] stage4_col76;
    logic [6:0] stage4_col77;
    logic [7:0] stage4_col78;
    logic [6:0] stage4_col79;
    logic [7:0] stage4_col80;
    logic [6:0] stage4_col81;
    logic [7:0] stage4_col82;
    logic [6:0] stage4_col83;
    logic [7:0] stage4_col84;
    logic [6:0] stage4_col85;
    logic [7:0] stage4_col86;
    logic [6:0] stage4_col87;
    logic [7:0] stage4_col88;
    logic [6:0] stage4_col89;
    logic [7:0] stage4_col90;
    logic [6:0] stage4_col91;
    logic [7:0] stage4_col92;
    logic [6:0] stage4_col93;
    logic [7:0] stage4_col94;
    logic [6:0] stage4_col95;
    logic [7:0] stage4_col96;
    logic [6:0] stage4_col97;
    logic [7:0] stage4_col98;
    logic [6:0] stage4_col99;
    logic [7:0] stage4_col100;
    logic [6:0] stage4_col101;
    logic [7:0] stage4_col102;
    logic [6:0] stage4_col103;
    logic [7:0] stage4_col104;
    logic [6:0] stage4_col105;
    logic [7:0] stage4_col106;
    logic [6:0] stage4_col107;
    logic [7:0] stage4_col108;
    logic [6:0] stage4_col109;
    logic [7:0] stage4_col110;
    logic [6:0] stage4_col111;
    logic [7:0] stage4_col112;
    logic [6:0] stage4_col113;
    logic [7:0] stage4_col114;
    logic [6:0] stage4_col115;
    logic [7:0] stage4_col116;
    logic [6:0] stage4_col117;
    logic [7:0] stage4_col118;
    logic [6:0] stage4_col119;
    logic [7:0] stage4_col120;
    logic [6:0] stage4_col121;
    logic [7:0] stage4_col122;
    logic [6:0] stage4_col123;
    logic [7:0] stage4_col124;
    logic [6:0] stage4_col125;
    logic [7:0] stage4_col126;
    logic [56:0] stage4_col127;

    // Stage 5 signals
    logic [0:0] stage5_col0;
    logic [0:0] stage5_col1;
    logic [0:0] stage5_col2;
    logic [0:0] stage5_col3;
    logic [0:0] stage5_col4;
    logic [1:0] stage5_col5;
    logic [0:0] stage5_col6;
    logic [2:0] stage5_col7;
    logic [1:0] stage5_col8;
    logic [1:0] stage5_col9;
    logic [1:0] stage5_col10;
    logic [1:0] stage5_col11;
    logic [1:0] stage5_col12;
    logic [1:0] stage5_col13;
    logic [1:0] stage5_col14;
    logic [1:0] stage5_col15;
    logic [1:0] stage5_col16;
    logic [1:0] stage5_col17;
    logic [1:0] stage5_col18;
    logic [1:0] stage5_col19;
    logic [1:0] stage5_col20;
    logic [1:0] stage5_col21;
    logic [1:0] stage5_col22;
    logic [1:0] stage5_col23;
    logic [1:0] stage5_col24;
    logic [1:0] stage5_col25;
    logic [1:0] stage5_col26;
    logic [1:0] stage5_col27;
    logic [3:0] stage5_col28;
    logic [2:0] stage5_col29;
    logic [2:0] stage5_col30;
    logic [2:0] stage5_col31;
    logic [2:0] stage5_col32;
    logic [2:0] stage5_col33;
    logic [2:0] stage5_col34;
    logic [2:0] stage5_col35;
    logic [2:0] stage5_col36;
    logic [2:0] stage5_col37;
    logic [2:0] stage5_col38;
    logic [2:0] stage5_col39;
    logic [2:0] stage5_col40;
    logic [4:0] stage5_col41;
    logic [3:0] stage5_col42;
    logic [3:0] stage5_col43;
    logic [3:0] stage5_col44;
    logic [3:0] stage5_col45;
    logic [3:0] stage5_col46;
    logic [3:0] stage5_col47;
    logic [3:0] stage5_col48;
    logic [3:0] stage5_col49;
    logic [3:0] stage5_col50;
    logic [3:0] stage5_col51;
    logic [3:0] stage5_col52;
    logic [3:0] stage5_col53;
    logic [3:0] stage5_col54;
    logic [3:0] stage5_col55;
    logic [3:0] stage5_col56;
    logic [3:0] stage5_col57;
    logic [3:0] stage5_col58;
    logic [5:0] stage5_col59;
    logic [4:0] stage5_col60;
    logic [4:0] stage5_col61;
    logic [4:0] stage5_col62;
    logic [4:0] stage5_col63;
    logic [5:0] stage5_col64;
    logic [4:0] stage5_col65;
    logic [5:0] stage5_col66;
    logic [4:0] stage5_col67;
    logic [5:0] stage5_col68;
    logic [4:0] stage5_col69;
    logic [5:0] stage5_col70;
    logic [4:0] stage5_col71;
    logic [5:0] stage5_col72;
    logic [4:0] stage5_col73;
    logic [5:0] stage5_col74;
    logic [4:0] stage5_col75;
    logic [5:0] stage5_col76;
    logic [4:0] stage5_col77;
    logic [5:0] stage5_col78;
    logic [4:0] stage5_col79;
    logic [5:0] stage5_col80;
    logic [4:0] stage5_col81;
    logic [5:0] stage5_col82;
    logic [4:0] stage5_col83;
    logic [5:0] stage5_col84;
    logic [4:0] stage5_col85;
    logic [5:0] stage5_col86;
    logic [4:0] stage5_col87;
    logic [5:0] stage5_col88;
    logic [4:0] stage5_col89;
    logic [5:0] stage5_col90;
    logic [4:0] stage5_col91;
    logic [5:0] stage5_col92;
    logic [4:0] stage5_col93;
    logic [5:0] stage5_col94;
    logic [4:0] stage5_col95;
    logic [5:0] stage5_col96;
    logic [4:0] stage5_col97;
    logic [5:0] stage5_col98;
    logic [4:0] stage5_col99;
    logic [5:0] stage5_col100;
    logic [4:0] stage5_col101;
    logic [5:0] stage5_col102;
    logic [4:0] stage5_col103;
    logic [5:0] stage5_col104;
    logic [4:0] stage5_col105;
    logic [5:0] stage5_col106;
    logic [4:0] stage5_col107;
    logic [5:0] stage5_col108;
    logic [4:0] stage5_col109;
    logic [5:0] stage5_col110;
    logic [4:0] stage5_col111;
    logic [5:0] stage5_col112;
    logic [4:0] stage5_col113;
    logic [5:0] stage5_col114;
    logic [4:0] stage5_col115;
    logic [5:0] stage5_col116;
    logic [4:0] stage5_col117;
    logic [5:0] stage5_col118;
    logic [4:0] stage5_col119;
    logic [5:0] stage5_col120;
    logic [4:0] stage5_col121;
    logic [5:0] stage5_col122;
    logic [4:0] stage5_col123;
    logic [5:0] stage5_col124;
    logic [4:0] stage5_col125;
    logic [5:0] stage5_col126;
    logic [58:0] stage5_col127;

    // Stage 6 signals
    logic [0:0] stage6_col0;
    logic [0:0] stage6_col1;
    logic [0:0] stage6_col2;
    logic [0:0] stage6_col3;
    logic [0:0] stage6_col4;
    logic [0:0] stage6_col5;
    logic [1:0] stage6_col6;
    logic [0:0] stage6_col7;
    logic [2:0] stage6_col8;
    logic [1:0] stage6_col9;
    logic [1:0] stage6_col10;
    logic [1:0] stage6_col11;
    logic [1:0] stage6_col12;
    logic [1:0] stage6_col13;
    logic [1:0] stage6_col14;
    logic [1:0] stage6_col15;
    logic [1:0] stage6_col16;
    logic [1:0] stage6_col17;
    logic [1:0] stage6_col18;
    logic [1:0] stage6_col19;
    logic [1:0] stage6_col20;
    logic [1:0] stage6_col21;
    logic [1:0] stage6_col22;
    logic [1:0] stage6_col23;
    logic [1:0] stage6_col24;
    logic [1:0] stage6_col25;
    logic [1:0] stage6_col26;
    logic [1:0] stage6_col27;
    logic [1:0] stage6_col28;
    logic [1:0] stage6_col29;
    logic [1:0] stage6_col30;
    logic [1:0] stage6_col31;
    logic [1:0] stage6_col32;
    logic [1:0] stage6_col33;
    logic [1:0] stage6_col34;
    logic [1:0] stage6_col35;
    logic [1:0] stage6_col36;
    logic [1:0] stage6_col37;
    logic [1:0] stage6_col38;
    logic [1:0] stage6_col39;
    logic [1:0] stage6_col40;
    logic [3:0] stage6_col41;
    logic [2:0] stage6_col42;
    logic [2:0] stage6_col43;
    logic [2:0] stage6_col44;
    logic [2:0] stage6_col45;
    logic [2:0] stage6_col46;
    logic [2:0] stage6_col47;
    logic [2:0] stage6_col48;
    logic [2:0] stage6_col49;
    logic [2:0] stage6_col50;
    logic [2:0] stage6_col51;
    logic [2:0] stage6_col52;
    logic [2:0] stage6_col53;
    logic [2:0] stage6_col54;
    logic [2:0] stage6_col55;
    logic [2:0] stage6_col56;
    logic [2:0] stage6_col57;
    logic [2:0] stage6_col58;
    logic [2:0] stage6_col59;
    logic [3:0] stage6_col60;
    logic [3:0] stage6_col61;
    logic [3:0] stage6_col62;
    logic [3:0] stage6_col63;
    logic [3:0] stage6_col64;
    logic [3:0] stage6_col65;
    logic [3:0] stage6_col66;
    logic [3:0] stage6_col67;
    logic [3:0] stage6_col68;
    logic [3:0] stage6_col69;
    logic [3:0] stage6_col70;
    logic [3:0] stage6_col71;
    logic [3:0] stage6_col72;
    logic [3:0] stage6_col73;
    logic [3:0] stage6_col74;
    logic [3:0] stage6_col75;
    logic [3:0] stage6_col76;
    logic [3:0] stage6_col77;
    logic [3:0] stage6_col78;
    logic [3:0] stage6_col79;
    logic [3:0] stage6_col80;
    logic [3:0] stage6_col81;
    logic [3:0] stage6_col82;
    logic [3:0] stage6_col83;
    logic [3:0] stage6_col84;
    logic [3:0] stage6_col85;
    logic [3:0] stage6_col86;
    logic [3:0] stage6_col87;
    logic [3:0] stage6_col88;
    logic [3:0] stage6_col89;
    logic [3:0] stage6_col90;
    logic [3:0] stage6_col91;
    logic [3:0] stage6_col92;
    logic [3:0] stage6_col93;
    logic [3:0] stage6_col94;
    logic [3:0] stage6_col95;
    logic [3:0] stage6_col96;
    logic [3:0] stage6_col97;
    logic [3:0] stage6_col98;
    logic [3:0] stage6_col99;
    logic [3:0] stage6_col100;
    logic [3:0] stage6_col101;
    logic [3:0] stage6_col102;
    logic [3:0] stage6_col103;
    logic [3:0] stage6_col104;
    logic [3:0] stage6_col105;
    logic [3:0] stage6_col106;
    logic [3:0] stage6_col107;
    logic [3:0] stage6_col108;
    logic [3:0] stage6_col109;
    logic [3:0] stage6_col110;
    logic [3:0] stage6_col111;
    logic [3:0] stage6_col112;
    logic [3:0] stage6_col113;
    logic [3:0] stage6_col114;
    logic [3:0] stage6_col115;
    logic [3:0] stage6_col116;
    logic [3:0] stage6_col117;
    logic [3:0] stage6_col118;
    logic [3:0] stage6_col119;
    logic [3:0] stage6_col120;
    logic [3:0] stage6_col121;
    logic [3:0] stage6_col122;
    logic [3:0] stage6_col123;
    logic [3:0] stage6_col124;
    logic [3:0] stage6_col125;
    logic [3:0] stage6_col126;
    logic [60:0] stage6_col127;

    // Stage 7 signals
    logic [0:0] stage7_col0;
    logic [0:0] stage7_col1;
    logic [0:0] stage7_col2;
    logic [0:0] stage7_col3;
    logic [0:0] stage7_col4;
    logic [0:0] stage7_col5;
    logic [0:0] stage7_col6;
    logic [1:0] stage7_col7;
    logic [0:0] stage7_col8;
    logic [2:0] stage7_col9;
    logic [1:0] stage7_col10;
    logic [1:0] stage7_col11;
    logic [1:0] stage7_col12;
    logic [1:0] stage7_col13;
    logic [1:0] stage7_col14;
    logic [1:0] stage7_col15;
    logic [1:0] stage7_col16;
    logic [1:0] stage7_col17;
    logic [1:0] stage7_col18;
    logic [1:0] stage7_col19;
    logic [1:0] stage7_col20;
    logic [1:0] stage7_col21;
    logic [1:0] stage7_col22;
    logic [1:0] stage7_col23;
    logic [1:0] stage7_col24;
    logic [1:0] stage7_col25;
    logic [1:0] stage7_col26;
    logic [1:0] stage7_col27;
    logic [1:0] stage7_col28;
    logic [1:0] stage7_col29;
    logic [1:0] stage7_col30;
    logic [1:0] stage7_col31;
    logic [1:0] stage7_col32;
    logic [1:0] stage7_col33;
    logic [1:0] stage7_col34;
    logic [1:0] stage7_col35;
    logic [1:0] stage7_col36;
    logic [1:0] stage7_col37;
    logic [1:0] stage7_col38;
    logic [1:0] stage7_col39;
    logic [1:0] stage7_col40;
    logic [1:0] stage7_col41;
    logic [1:0] stage7_col42;
    logic [1:0] stage7_col43;
    logic [1:0] stage7_col44;
    logic [1:0] stage7_col45;
    logic [1:0] stage7_col46;
    logic [1:0] stage7_col47;
    logic [1:0] stage7_col48;
    logic [1:0] stage7_col49;
    logic [1:0] stage7_col50;
    logic [1:0] stage7_col51;
    logic [1:0] stage7_col52;
    logic [1:0] stage7_col53;
    logic [1:0] stage7_col54;
    logic [1:0] stage7_col55;
    logic [1:0] stage7_col56;
    logic [1:0] stage7_col57;
    logic [1:0] stage7_col58;
    logic [1:0] stage7_col59;
    logic [2:0] stage7_col60;
    logic [2:0] stage7_col61;
    logic [2:0] stage7_col62;
    logic [2:0] stage7_col63;
    logic [2:0] stage7_col64;
    logic [2:0] stage7_col65;
    logic [2:0] stage7_col66;
    logic [2:0] stage7_col67;
    logic [2:0] stage7_col68;
    logic [2:0] stage7_col69;
    logic [2:0] stage7_col70;
    logic [2:0] stage7_col71;
    logic [2:0] stage7_col72;
    logic [2:0] stage7_col73;
    logic [2:0] stage7_col74;
    logic [2:0] stage7_col75;
    logic [2:0] stage7_col76;
    logic [2:0] stage7_col77;
    logic [2:0] stage7_col78;
    logic [2:0] stage7_col79;
    logic [2:0] stage7_col80;
    logic [2:0] stage7_col81;
    logic [2:0] stage7_col82;
    logic [2:0] stage7_col83;
    logic [2:0] stage7_col84;
    logic [2:0] stage7_col85;
    logic [2:0] stage7_col86;
    logic [2:0] stage7_col87;
    logic [2:0] stage7_col88;
    logic [2:0] stage7_col89;
    logic [2:0] stage7_col90;
    logic [2:0] stage7_col91;
    logic [2:0] stage7_col92;
    logic [2:0] stage7_col93;
    logic [2:0] stage7_col94;
    logic [2:0] stage7_col95;
    logic [2:0] stage7_col96;
    logic [2:0] stage7_col97;
    logic [2:0] stage7_col98;
    logic [2:0] stage7_col99;
    logic [2:0] stage7_col100;
    logic [2:0] stage7_col101;
    logic [2:0] stage7_col102;
    logic [2:0] stage7_col103;
    logic [2:0] stage7_col104;
    logic [2:0] stage7_col105;
    logic [2:0] stage7_col106;
    logic [2:0] stage7_col107;
    logic [2:0] stage7_col108;
    logic [2:0] stage7_col109;
    logic [2:0] stage7_col110;
    logic [2:0] stage7_col111;
    logic [2:0] stage7_col112;
    logic [2:0] stage7_col113;
    logic [2:0] stage7_col114;
    logic [2:0] stage7_col115;
    logic [2:0] stage7_col116;
    logic [2:0] stage7_col117;
    logic [2:0] stage7_col118;
    logic [2:0] stage7_col119;
    logic [2:0] stage7_col120;
    logic [2:0] stage7_col121;
    logic [2:0] stage7_col122;
    logic [2:0] stage7_col123;
    logic [2:0] stage7_col124;
    logic [2:0] stage7_col125;
    logic [2:0] stage7_col126;
    logic [61:0] stage7_col127;

    // Stage 8 signals
    logic [0:0] stage8_col0;
    logic [0:0] stage8_col1;
    logic [0:0] stage8_col2;
    logic [0:0] stage8_col3;
    logic [0:0] stage8_col4;
    logic [0:0] stage8_col5;
    logic [0:0] stage8_col6;
    logic [0:0] stage8_col7;
    logic [1:0] stage8_col8;
    logic [0:0] stage8_col9;
    logic [1:0] stage8_col10;
    logic [1:0] stage8_col11;
    logic [1:0] stage8_col12;
    logic [1:0] stage8_col13;
    logic [1:0] stage8_col14;
    logic [1:0] stage8_col15;
    logic [1:0] stage8_col16;
    logic [1:0] stage8_col17;
    logic [1:0] stage8_col18;
    logic [1:0] stage8_col19;
    logic [1:0] stage8_col20;
    logic [1:0] stage8_col21;
    logic [1:0] stage8_col22;
    logic [1:0] stage8_col23;
    logic [1:0] stage8_col24;
    logic [1:0] stage8_col25;
    logic [1:0] stage8_col26;
    logic [1:0] stage8_col27;
    logic [1:0] stage8_col28;
    logic [1:0] stage8_col29;
    logic [1:0] stage8_col30;
    logic [1:0] stage8_col31;
    logic [1:0] stage8_col32;
    logic [1:0] stage8_col33;
    logic [1:0] stage8_col34;
    logic [1:0] stage8_col35;
    logic [1:0] stage8_col36;
    logic [1:0] stage8_col37;
    logic [1:0] stage8_col38;
    logic [1:0] stage8_col39;
    logic [1:0] stage8_col40;
    logic [1:0] stage8_col41;
    logic [1:0] stage8_col42;
    logic [1:0] stage8_col43;
    logic [1:0] stage8_col44;
    logic [1:0] stage8_col45;
    logic [1:0] stage8_col46;
    logic [1:0] stage8_col47;
    logic [1:0] stage8_col48;
    logic [1:0] stage8_col49;
    logic [1:0] stage8_col50;
    logic [1:0] stage8_col51;
    logic [1:0] stage8_col52;
    logic [1:0] stage8_col53;
    logic [1:0] stage8_col54;
    logic [1:0] stage8_col55;
    logic [1:0] stage8_col56;
    logic [1:0] stage8_col57;
    logic [1:0] stage8_col58;
    logic [1:0] stage8_col59;
    logic [1:0] stage8_col60;
    logic [1:0] stage8_col61;
    logic [1:0] stage8_col62;
    logic [1:0] stage8_col63;
    logic [1:0] stage8_col64;
    logic [1:0] stage8_col65;
    logic [1:0] stage8_col66;
    logic [1:0] stage8_col67;
    logic [1:0] stage8_col68;
    logic [1:0] stage8_col69;
    logic [1:0] stage8_col70;
    logic [1:0] stage8_col71;
    logic [1:0] stage8_col72;
    logic [1:0] stage8_col73;
    logic [1:0] stage8_col74;
    logic [1:0] stage8_col75;
    logic [1:0] stage8_col76;
    logic [1:0] stage8_col77;
    logic [1:0] stage8_col78;
    logic [1:0] stage8_col79;
    logic [1:0] stage8_col80;
    logic [1:0] stage8_col81;
    logic [1:0] stage8_col82;
    logic [1:0] stage8_col83;
    logic [1:0] stage8_col84;
    logic [1:0] stage8_col85;
    logic [1:0] stage8_col86;
    logic [1:0] stage8_col87;
    logic [1:0] stage8_col88;
    logic [1:0] stage8_col89;
    logic [1:0] stage8_col90;
    logic [1:0] stage8_col91;
    logic [1:0] stage8_col92;
    logic [1:0] stage8_col93;
    logic [1:0] stage8_col94;
    logic [1:0] stage8_col95;
    logic [1:0] stage8_col96;
    logic [1:0] stage8_col97;
    logic [1:0] stage8_col98;
    logic [1:0] stage8_col99;
    logic [1:0] stage8_col100;
    logic [1:0] stage8_col101;
    logic [1:0] stage8_col102;
    logic [1:0] stage8_col103;
    logic [1:0] stage8_col104;
    logic [1:0] stage8_col105;
    logic [1:0] stage8_col106;
    logic [1:0] stage8_col107;
    logic [1:0] stage8_col108;
    logic [1:0] stage8_col109;
    logic [1:0] stage8_col110;
    logic [1:0] stage8_col111;
    logic [1:0] stage8_col112;
    logic [1:0] stage8_col113;
    logic [1:0] stage8_col114;
    logic [1:0] stage8_col115;
    logic [1:0] stage8_col116;
    logic [1:0] stage8_col117;
    logic [1:0] stage8_col118;
    logic [1:0] stage8_col119;
    logic [1:0] stage8_col120;
    logic [1:0] stage8_col121;
    logic [1:0] stage8_col122;
    logic [1:0] stage8_col123;
    logic [1:0] stage8_col124;
    logic [1:0] stage8_col125;
    logic [1:0] stage8_col126;
    logic [62:0] stage8_col127;

    // Stage 0: Partial Product Assignment
    // Combinational assignment
    always_comb begin
        stage0_col0[0] = cpl[0];
        stage0_col0[1] = pp[0][0];
        stage0_col1[0] = pp[0][1];
        stage0_col2[0] = pp[0][2];
        stage0_col2[1] = cpl[1];
        stage0_col2[2] = pp[1][0];
        stage0_col3[0] = pp[0][3];
        stage0_col3[1] = pp[1][1];
        stage0_col4[0] = pp[0][4];
        stage0_col4[1] = pp[1][2];
        stage0_col4[2] = cpl[2];
        stage0_col4[3] = pp[2][0];
        stage0_col5[0] = pp[0][5];
        stage0_col5[1] = pp[1][3];
        stage0_col5[2] = pp[2][1];
        stage0_col6[0] = pp[0][6];
        stage0_col6[1] = pp[1][4];
        stage0_col6[2] = pp[2][2];
        stage0_col6[3] = cpl[3];
        stage0_col6[4] = pp[3][0];
        stage0_col7[0] = pp[0][7];
        stage0_col7[1] = pp[1][5];
        stage0_col7[2] = pp[2][3];
        stage0_col7[3] = pp[3][1];
        stage0_col8[0] = pp[0][8];
        stage0_col8[1] = pp[1][6];
        stage0_col8[2] = pp[2][4];
        stage0_col8[3] = pp[3][2];
        stage0_col8[4] = cpl[4];
        stage0_col8[5] = pp[4][0];
        stage0_col9[0] = pp[0][9];
        stage0_col9[1] = pp[1][7];
        stage0_col9[2] = pp[2][5];
        stage0_col9[3] = pp[3][3];
        stage0_col9[4] = pp[4][1];
        stage0_col10[0] = pp[0][10];
        stage0_col10[1] = pp[1][8];
        stage0_col10[2] = pp[2][6];
        stage0_col10[3] = pp[3][4];
        stage0_col10[4] = pp[4][2];
        stage0_col10[5] = cpl[5];
        stage0_col10[6] = pp[5][0];
        stage0_col11[0] = pp[0][11];
        stage0_col11[1] = pp[1][9];
        stage0_col11[2] = pp[2][7];
        stage0_col11[3] = pp[3][5];
        stage0_col11[4] = pp[4][3];
        stage0_col11[5] = pp[5][1];
        stage0_col12[0] = pp[0][12];
        stage0_col12[1] = pp[1][10];
        stage0_col12[2] = pp[2][8];
        stage0_col12[3] = pp[3][6];
        stage0_col12[4] = pp[4][4];
        stage0_col12[5] = pp[5][2];
        stage0_col12[6] = cpl[6];
        stage0_col12[7] = pp[6][0];
        stage0_col13[0] = pp[0][13];
        stage0_col13[1] = pp[1][11];
        stage0_col13[2] = pp[2][9];
        stage0_col13[3] = pp[3][7];
        stage0_col13[4] = pp[4][5];
        stage0_col13[5] = pp[5][3];
        stage0_col13[6] = pp[6][1];
        stage0_col14[0] = pp[0][14];
        stage0_col14[1] = pp[1][12];
        stage0_col14[2] = pp[2][10];
        stage0_col14[3] = pp[3][8];
        stage0_col14[4] = pp[4][6];
        stage0_col14[5] = pp[5][4];
        stage0_col14[6] = pp[6][2];
        stage0_col14[7] = cpl[7];
        stage0_col14[8] = pp[7][0];
        stage0_col15[0] = pp[0][15];
        stage0_col15[1] = pp[1][13];
        stage0_col15[2] = pp[2][11];
        stage0_col15[3] = pp[3][9];
        stage0_col15[4] = pp[4][7];
        stage0_col15[5] = pp[5][5];
        stage0_col15[6] = pp[6][3];
        stage0_col15[7] = pp[7][1];
        stage0_col16[0] = pp[0][16];
        stage0_col16[1] = pp[1][14];
        stage0_col16[2] = pp[2][12];
        stage0_col16[3] = pp[3][10];
        stage0_col16[4] = pp[4][8];
        stage0_col16[5] = pp[5][6];
        stage0_col16[6] = pp[6][4];
        stage0_col16[7] = pp[7][2];
        stage0_col16[8] = cpl[8];
        stage0_col16[9] = pp[8][0];
        stage0_col17[0] = pp[0][17];
        stage0_col17[1] = pp[1][15];
        stage0_col17[2] = pp[2][13];
        stage0_col17[3] = pp[3][11];
        stage0_col17[4] = pp[4][9];
        stage0_col17[5] = pp[5][7];
        stage0_col17[6] = pp[6][5];
        stage0_col17[7] = pp[7][3];
        stage0_col17[8] = pp[8][1];
        stage0_col18[0] = pp[0][18];
        stage0_col18[1] = pp[1][16];
        stage0_col18[2] = pp[2][14];
        stage0_col18[3] = pp[3][12];
        stage0_col18[4] = pp[4][10];
        stage0_col18[5] = pp[5][8];
        stage0_col18[6] = pp[6][6];
        stage0_col18[7] = pp[7][4];
        stage0_col18[8] = pp[8][2];
        stage0_col18[9] = cpl[9];
        stage0_col18[10] = pp[9][0];
        stage0_col19[0] = pp[0][19];
        stage0_col19[1] = pp[1][17];
        stage0_col19[2] = pp[2][15];
        stage0_col19[3] = pp[3][13];
        stage0_col19[4] = pp[4][11];
        stage0_col19[5] = pp[5][9];
        stage0_col19[6] = pp[6][7];
        stage0_col19[7] = pp[7][5];
        stage0_col19[8] = pp[8][3];
        stage0_col19[9] = pp[9][1];
        stage0_col20[0] = pp[0][20];
        stage0_col20[1] = pp[1][18];
        stage0_col20[2] = pp[2][16];
        stage0_col20[3] = pp[3][14];
        stage0_col20[4] = pp[4][12];
        stage0_col20[5] = pp[5][10];
        stage0_col20[6] = pp[6][8];
        stage0_col20[7] = pp[7][6];
        stage0_col20[8] = pp[8][4];
        stage0_col20[9] = pp[9][2];
        stage0_col20[10] = cpl[10];
        stage0_col20[11] = pp[10][0];
        stage0_col21[0] = pp[0][21];
        stage0_col21[1] = pp[1][19];
        stage0_col21[2] = pp[2][17];
        stage0_col21[3] = pp[3][15];
        stage0_col21[4] = pp[4][13];
        stage0_col21[5] = pp[5][11];
        stage0_col21[6] = pp[6][9];
        stage0_col21[7] = pp[7][7];
        stage0_col21[8] = pp[8][5];
        stage0_col21[9] = pp[9][3];
        stage0_col21[10] = pp[10][1];
        stage0_col22[0] = pp[0][22];
        stage0_col22[1] = pp[1][20];
        stage0_col22[2] = pp[2][18];
        stage0_col22[3] = pp[3][16];
        stage0_col22[4] = pp[4][14];
        stage0_col22[5] = pp[5][12];
        stage0_col22[6] = pp[6][10];
        stage0_col22[7] = pp[7][8];
        stage0_col22[8] = pp[8][6];
        stage0_col22[9] = pp[9][4];
        stage0_col22[10] = pp[10][2];
        stage0_col22[11] = cpl[11];
        stage0_col22[12] = pp[11][0];
        stage0_col23[0] = pp[0][23];
        stage0_col23[1] = pp[1][21];
        stage0_col23[2] = pp[2][19];
        stage0_col23[3] = pp[3][17];
        stage0_col23[4] = pp[4][15];
        stage0_col23[5] = pp[5][13];
        stage0_col23[6] = pp[6][11];
        stage0_col23[7] = pp[7][9];
        stage0_col23[8] = pp[8][7];
        stage0_col23[9] = pp[9][5];
        stage0_col23[10] = pp[10][3];
        stage0_col23[11] = pp[11][1];
        stage0_col24[0] = pp[0][24];
        stage0_col24[1] = pp[1][22];
        stage0_col24[2] = pp[2][20];
        stage0_col24[3] = pp[3][18];
        stage0_col24[4] = pp[4][16];
        stage0_col24[5] = pp[5][14];
        stage0_col24[6] = pp[6][12];
        stage0_col24[7] = pp[7][10];
        stage0_col24[8] = pp[8][8];
        stage0_col24[9] = pp[9][6];
        stage0_col24[10] = pp[10][4];
        stage0_col24[11] = pp[11][2];
        stage0_col24[12] = cpl[12];
        stage0_col24[13] = pp[12][0];
        stage0_col25[0] = pp[0][25];
        stage0_col25[1] = pp[1][23];
        stage0_col25[2] = pp[2][21];
        stage0_col25[3] = pp[3][19];
        stage0_col25[4] = pp[4][17];
        stage0_col25[5] = pp[5][15];
        stage0_col25[6] = pp[6][13];
        stage0_col25[7] = pp[7][11];
        stage0_col25[8] = pp[8][9];
        stage0_col25[9] = pp[9][7];
        stage0_col25[10] = pp[10][5];
        stage0_col25[11] = pp[11][3];
        stage0_col25[12] = pp[12][1];
        stage0_col26[0] = pp[0][26];
        stage0_col26[1] = pp[1][24];
        stage0_col26[2] = pp[2][22];
        stage0_col26[3] = pp[3][20];
        stage0_col26[4] = pp[4][18];
        stage0_col26[5] = pp[5][16];
        stage0_col26[6] = pp[6][14];
        stage0_col26[7] = pp[7][12];
        stage0_col26[8] = pp[8][10];
        stage0_col26[9] = pp[9][8];
        stage0_col26[10] = pp[10][6];
        stage0_col26[11] = pp[11][4];
        stage0_col26[12] = pp[12][2];
        stage0_col26[13] = cpl[13];
        stage0_col26[14] = pp[13][0];
        stage0_col27[0] = pp[0][27];
        stage0_col27[1] = pp[1][25];
        stage0_col27[2] = pp[2][23];
        stage0_col27[3] = pp[3][21];
        stage0_col27[4] = pp[4][19];
        stage0_col27[5] = pp[5][17];
        stage0_col27[6] = pp[6][15];
        stage0_col27[7] = pp[7][13];
        stage0_col27[8] = pp[8][11];
        stage0_col27[9] = pp[9][9];
        stage0_col27[10] = pp[10][7];
        stage0_col27[11] = pp[11][5];
        stage0_col27[12] = pp[12][3];
        stage0_col27[13] = pp[13][1];
        stage0_col28[0] = pp[0][28];
        stage0_col28[1] = pp[1][26];
        stage0_col28[2] = pp[2][24];
        stage0_col28[3] = pp[3][22];
        stage0_col28[4] = pp[4][20];
        stage0_col28[5] = pp[5][18];
        stage0_col28[6] = pp[6][16];
        stage0_col28[7] = pp[7][14];
        stage0_col28[8] = pp[8][12];
        stage0_col28[9] = pp[9][10];
        stage0_col28[10] = pp[10][8];
        stage0_col28[11] = pp[11][6];
        stage0_col28[12] = pp[12][4];
        stage0_col28[13] = pp[13][2];
        stage0_col28[14] = cpl[14];
        stage0_col28[15] = pp[14][0];
        stage0_col29[0] = pp[0][29];
        stage0_col29[1] = pp[1][27];
        stage0_col29[2] = pp[2][25];
        stage0_col29[3] = pp[3][23];
        stage0_col29[4] = pp[4][21];
        stage0_col29[5] = pp[5][19];
        stage0_col29[6] = pp[6][17];
        stage0_col29[7] = pp[7][15];
        stage0_col29[8] = pp[8][13];
        stage0_col29[9] = pp[9][11];
        stage0_col29[10] = pp[10][9];
        stage0_col29[11] = pp[11][7];
        stage0_col29[12] = pp[12][5];
        stage0_col29[13] = pp[13][3];
        stage0_col29[14] = pp[14][1];
        stage0_col30[0] = pp[0][30];
        stage0_col30[1] = pp[1][28];
        stage0_col30[2] = pp[2][26];
        stage0_col30[3] = pp[3][24];
        stage0_col30[4] = pp[4][22];
        stage0_col30[5] = pp[5][20];
        stage0_col30[6] = pp[6][18];
        stage0_col30[7] = pp[7][16];
        stage0_col30[8] = pp[8][14];
        stage0_col30[9] = pp[9][12];
        stage0_col30[10] = pp[10][10];
        stage0_col30[11] = pp[11][8];
        stage0_col30[12] = pp[12][6];
        stage0_col30[13] = pp[13][4];
        stage0_col30[14] = pp[14][2];
        stage0_col30[15] = cpl[15];
        stage0_col30[16] = pp[15][0];
        stage0_col31[0] = pp[0][31];
        stage0_col31[1] = pp[1][29];
        stage0_col31[2] = pp[2][27];
        stage0_col31[3] = pp[3][25];
        stage0_col31[4] = pp[4][23];
        stage0_col31[5] = pp[5][21];
        stage0_col31[6] = pp[6][19];
        stage0_col31[7] = pp[7][17];
        stage0_col31[8] = pp[8][15];
        stage0_col31[9] = pp[9][13];
        stage0_col31[10] = pp[10][11];
        stage0_col31[11] = pp[11][9];
        stage0_col31[12] = pp[12][7];
        stage0_col31[13] = pp[13][5];
        stage0_col31[14] = pp[14][3];
        stage0_col31[15] = pp[15][1];
        stage0_col32[0] = pp[0][32];
        stage0_col32[1] = pp[1][30];
        stage0_col32[2] = pp[2][28];
        stage0_col32[3] = pp[3][26];
        stage0_col32[4] = pp[4][24];
        stage0_col32[5] = pp[5][22];
        stage0_col32[6] = pp[6][20];
        stage0_col32[7] = pp[7][18];
        stage0_col32[8] = pp[8][16];
        stage0_col32[9] = pp[9][14];
        stage0_col32[10] = pp[10][12];
        stage0_col32[11] = pp[11][10];
        stage0_col32[12] = pp[12][8];
        stage0_col32[13] = pp[13][6];
        stage0_col32[14] = pp[14][4];
        stage0_col32[15] = pp[15][2];
        stage0_col32[16] = cpl[16];
        stage0_col32[17] = pp[16][0];
        stage0_col33[0] = pp[0][33];
        stage0_col33[1] = pp[1][31];
        stage0_col33[2] = pp[2][29];
        stage0_col33[3] = pp[3][27];
        stage0_col33[4] = pp[4][25];
        stage0_col33[5] = pp[5][23];
        stage0_col33[6] = pp[6][21];
        stage0_col33[7] = pp[7][19];
        stage0_col33[8] = pp[8][17];
        stage0_col33[9] = pp[9][15];
        stage0_col33[10] = pp[10][13];
        stage0_col33[11] = pp[11][11];
        stage0_col33[12] = pp[12][9];
        stage0_col33[13] = pp[13][7];
        stage0_col33[14] = pp[14][5];
        stage0_col33[15] = pp[15][3];
        stage0_col33[16] = pp[16][1];
        stage0_col34[0] = pp[0][34];
        stage0_col34[1] = pp[1][32];
        stage0_col34[2] = pp[2][30];
        stage0_col34[3] = pp[3][28];
        stage0_col34[4] = pp[4][26];
        stage0_col34[5] = pp[5][24];
        stage0_col34[6] = pp[6][22];
        stage0_col34[7] = pp[7][20];
        stage0_col34[8] = pp[8][18];
        stage0_col34[9] = pp[9][16];
        stage0_col34[10] = pp[10][14];
        stage0_col34[11] = pp[11][12];
        stage0_col34[12] = pp[12][10];
        stage0_col34[13] = pp[13][8];
        stage0_col34[14] = pp[14][6];
        stage0_col34[15] = pp[15][4];
        stage0_col34[16] = pp[16][2];
        stage0_col34[17] = cpl[17];
        stage0_col34[18] = pp[17][0];
        stage0_col35[0] = pp[0][35];
        stage0_col35[1] = pp[1][33];
        stage0_col35[2] = pp[2][31];
        stage0_col35[3] = pp[3][29];
        stage0_col35[4] = pp[4][27];
        stage0_col35[5] = pp[5][25];
        stage0_col35[6] = pp[6][23];
        stage0_col35[7] = pp[7][21];
        stage0_col35[8] = pp[8][19];
        stage0_col35[9] = pp[9][17];
        stage0_col35[10] = pp[10][15];
        stage0_col35[11] = pp[11][13];
        stage0_col35[12] = pp[12][11];
        stage0_col35[13] = pp[13][9];
        stage0_col35[14] = pp[14][7];
        stage0_col35[15] = pp[15][5];
        stage0_col35[16] = pp[16][3];
        stage0_col35[17] = pp[17][1];
        stage0_col36[0] = pp[0][36];
        stage0_col36[1] = pp[1][34];
        stage0_col36[2] = pp[2][32];
        stage0_col36[3] = pp[3][30];
        stage0_col36[4] = pp[4][28];
        stage0_col36[5] = pp[5][26];
        stage0_col36[6] = pp[6][24];
        stage0_col36[7] = pp[7][22];
        stage0_col36[8] = pp[8][20];
        stage0_col36[9] = pp[9][18];
        stage0_col36[10] = pp[10][16];
        stage0_col36[11] = pp[11][14];
        stage0_col36[12] = pp[12][12];
        stage0_col36[13] = pp[13][10];
        stage0_col36[14] = pp[14][8];
        stage0_col36[15] = pp[15][6];
        stage0_col36[16] = pp[16][4];
        stage0_col36[17] = pp[17][2];
        stage0_col36[18] = cpl[18];
        stage0_col36[19] = pp[18][0];
        stage0_col37[0] = pp[0][37];
        stage0_col37[1] = pp[1][35];
        stage0_col37[2] = pp[2][33];
        stage0_col37[3] = pp[3][31];
        stage0_col37[4] = pp[4][29];
        stage0_col37[5] = pp[5][27];
        stage0_col37[6] = pp[6][25];
        stage0_col37[7] = pp[7][23];
        stage0_col37[8] = pp[8][21];
        stage0_col37[9] = pp[9][19];
        stage0_col37[10] = pp[10][17];
        stage0_col37[11] = pp[11][15];
        stage0_col37[12] = pp[12][13];
        stage0_col37[13] = pp[13][11];
        stage0_col37[14] = pp[14][9];
        stage0_col37[15] = pp[15][7];
        stage0_col37[16] = pp[16][5];
        stage0_col37[17] = pp[17][3];
        stage0_col37[18] = pp[18][1];
        stage0_col38[0] = pp[0][38];
        stage0_col38[1] = pp[1][36];
        stage0_col38[2] = pp[2][34];
        stage0_col38[3] = pp[3][32];
        stage0_col38[4] = pp[4][30];
        stage0_col38[5] = pp[5][28];
        stage0_col38[6] = pp[6][26];
        stage0_col38[7] = pp[7][24];
        stage0_col38[8] = pp[8][22];
        stage0_col38[9] = pp[9][20];
        stage0_col38[10] = pp[10][18];
        stage0_col38[11] = pp[11][16];
        stage0_col38[12] = pp[12][14];
        stage0_col38[13] = pp[13][12];
        stage0_col38[14] = pp[14][10];
        stage0_col38[15] = pp[15][8];
        stage0_col38[16] = pp[16][6];
        stage0_col38[17] = pp[17][4];
        stage0_col38[18] = pp[18][2];
        stage0_col38[19] = cpl[19];
        stage0_col38[20] = pp[19][0];
        stage0_col39[0] = pp[0][39];
        stage0_col39[1] = pp[1][37];
        stage0_col39[2] = pp[2][35];
        stage0_col39[3] = pp[3][33];
        stage0_col39[4] = pp[4][31];
        stage0_col39[5] = pp[5][29];
        stage0_col39[6] = pp[6][27];
        stage0_col39[7] = pp[7][25];
        stage0_col39[8] = pp[8][23];
        stage0_col39[9] = pp[9][21];
        stage0_col39[10] = pp[10][19];
        stage0_col39[11] = pp[11][17];
        stage0_col39[12] = pp[12][15];
        stage0_col39[13] = pp[13][13];
        stage0_col39[14] = pp[14][11];
        stage0_col39[15] = pp[15][9];
        stage0_col39[16] = pp[16][7];
        stage0_col39[17] = pp[17][5];
        stage0_col39[18] = pp[18][3];
        stage0_col39[19] = pp[19][1];
        stage0_col40[0] = pp[0][40];
        stage0_col40[1] = pp[1][38];
        stage0_col40[2] = pp[2][36];
        stage0_col40[3] = pp[3][34];
        stage0_col40[4] = pp[4][32];
        stage0_col40[5] = pp[5][30];
        stage0_col40[6] = pp[6][28];
        stage0_col40[7] = pp[7][26];
        stage0_col40[8] = pp[8][24];
        stage0_col40[9] = pp[9][22];
        stage0_col40[10] = pp[10][20];
        stage0_col40[11] = pp[11][18];
        stage0_col40[12] = pp[12][16];
        stage0_col40[13] = pp[13][14];
        stage0_col40[14] = pp[14][12];
        stage0_col40[15] = pp[15][10];
        stage0_col40[16] = pp[16][8];
        stage0_col40[17] = pp[17][6];
        stage0_col40[18] = pp[18][4];
        stage0_col40[19] = pp[19][2];
        stage0_col40[20] = cpl[20];
        stage0_col40[21] = pp[20][0];
        stage0_col41[0] = pp[0][41];
        stage0_col41[1] = pp[1][39];
        stage0_col41[2] = pp[2][37];
        stage0_col41[3] = pp[3][35];
        stage0_col41[4] = pp[4][33];
        stage0_col41[5] = pp[5][31];
        stage0_col41[6] = pp[6][29];
        stage0_col41[7] = pp[7][27];
        stage0_col41[8] = pp[8][25];
        stage0_col41[9] = pp[9][23];
        stage0_col41[10] = pp[10][21];
        stage0_col41[11] = pp[11][19];
        stage0_col41[12] = pp[12][17];
        stage0_col41[13] = pp[13][15];
        stage0_col41[14] = pp[14][13];
        stage0_col41[15] = pp[15][11];
        stage0_col41[16] = pp[16][9];
        stage0_col41[17] = pp[17][7];
        stage0_col41[18] = pp[18][5];
        stage0_col41[19] = pp[19][3];
        stage0_col41[20] = pp[20][1];
        stage0_col42[0] = pp[0][42];
        stage0_col42[1] = pp[1][40];
        stage0_col42[2] = pp[2][38];
        stage0_col42[3] = pp[3][36];
        stage0_col42[4] = pp[4][34];
        stage0_col42[5] = pp[5][32];
        stage0_col42[6] = pp[6][30];
        stage0_col42[7] = pp[7][28];
        stage0_col42[8] = pp[8][26];
        stage0_col42[9] = pp[9][24];
        stage0_col42[10] = pp[10][22];
        stage0_col42[11] = pp[11][20];
        stage0_col42[12] = pp[12][18];
        stage0_col42[13] = pp[13][16];
        stage0_col42[14] = pp[14][14];
        stage0_col42[15] = pp[15][12];
        stage0_col42[16] = pp[16][10];
        stage0_col42[17] = pp[17][8];
        stage0_col42[18] = pp[18][6];
        stage0_col42[19] = pp[19][4];
        stage0_col42[20] = pp[20][2];
        stage0_col42[21] = cpl[21];
        stage0_col42[22] = pp[21][0];
        stage0_col43[0] = pp[0][43];
        stage0_col43[1] = pp[1][41];
        stage0_col43[2] = pp[2][39];
        stage0_col43[3] = pp[3][37];
        stage0_col43[4] = pp[4][35];
        stage0_col43[5] = pp[5][33];
        stage0_col43[6] = pp[6][31];
        stage0_col43[7] = pp[7][29];
        stage0_col43[8] = pp[8][27];
        stage0_col43[9] = pp[9][25];
        stage0_col43[10] = pp[10][23];
        stage0_col43[11] = pp[11][21];
        stage0_col43[12] = pp[12][19];
        stage0_col43[13] = pp[13][17];
        stage0_col43[14] = pp[14][15];
        stage0_col43[15] = pp[15][13];
        stage0_col43[16] = pp[16][11];
        stage0_col43[17] = pp[17][9];
        stage0_col43[18] = pp[18][7];
        stage0_col43[19] = pp[19][5];
        stage0_col43[20] = pp[20][3];
        stage0_col43[21] = pp[21][1];
        stage0_col44[0] = pp[0][44];
        stage0_col44[1] = pp[1][42];
        stage0_col44[2] = pp[2][40];
        stage0_col44[3] = pp[3][38];
        stage0_col44[4] = pp[4][36];
        stage0_col44[5] = pp[5][34];
        stage0_col44[6] = pp[6][32];
        stage0_col44[7] = pp[7][30];
        stage0_col44[8] = pp[8][28];
        stage0_col44[9] = pp[9][26];
        stage0_col44[10] = pp[10][24];
        stage0_col44[11] = pp[11][22];
        stage0_col44[12] = pp[12][20];
        stage0_col44[13] = pp[13][18];
        stage0_col44[14] = pp[14][16];
        stage0_col44[15] = pp[15][14];
        stage0_col44[16] = pp[16][12];
        stage0_col44[17] = pp[17][10];
        stage0_col44[18] = pp[18][8];
        stage0_col44[19] = pp[19][6];
        stage0_col44[20] = pp[20][4];
        stage0_col44[21] = pp[21][2];
        stage0_col44[22] = cpl[22];
        stage0_col44[23] = pp[22][0];
        stage0_col45[0] = pp[0][45];
        stage0_col45[1] = pp[1][43];
        stage0_col45[2] = pp[2][41];
        stage0_col45[3] = pp[3][39];
        stage0_col45[4] = pp[4][37];
        stage0_col45[5] = pp[5][35];
        stage0_col45[6] = pp[6][33];
        stage0_col45[7] = pp[7][31];
        stage0_col45[8] = pp[8][29];
        stage0_col45[9] = pp[9][27];
        stage0_col45[10] = pp[10][25];
        stage0_col45[11] = pp[11][23];
        stage0_col45[12] = pp[12][21];
        stage0_col45[13] = pp[13][19];
        stage0_col45[14] = pp[14][17];
        stage0_col45[15] = pp[15][15];
        stage0_col45[16] = pp[16][13];
        stage0_col45[17] = pp[17][11];
        stage0_col45[18] = pp[18][9];
        stage0_col45[19] = pp[19][7];
        stage0_col45[20] = pp[20][5];
        stage0_col45[21] = pp[21][3];
        stage0_col45[22] = pp[22][1];
        stage0_col46[0] = pp[0][46];
        stage0_col46[1] = pp[1][44];
        stage0_col46[2] = pp[2][42];
        stage0_col46[3] = pp[3][40];
        stage0_col46[4] = pp[4][38];
        stage0_col46[5] = pp[5][36];
        stage0_col46[6] = pp[6][34];
        stage0_col46[7] = pp[7][32];
        stage0_col46[8] = pp[8][30];
        stage0_col46[9] = pp[9][28];
        stage0_col46[10] = pp[10][26];
        stage0_col46[11] = pp[11][24];
        stage0_col46[12] = pp[12][22];
        stage0_col46[13] = pp[13][20];
        stage0_col46[14] = pp[14][18];
        stage0_col46[15] = pp[15][16];
        stage0_col46[16] = pp[16][14];
        stage0_col46[17] = pp[17][12];
        stage0_col46[18] = pp[18][10];
        stage0_col46[19] = pp[19][8];
        stage0_col46[20] = pp[20][6];
        stage0_col46[21] = pp[21][4];
        stage0_col46[22] = pp[22][2];
        stage0_col46[23] = cpl[23];
        stage0_col46[24] = pp[23][0];
        stage0_col47[0] = pp[0][47];
        stage0_col47[1] = pp[1][45];
        stage0_col47[2] = pp[2][43];
        stage0_col47[3] = pp[3][41];
        stage0_col47[4] = pp[4][39];
        stage0_col47[5] = pp[5][37];
        stage0_col47[6] = pp[6][35];
        stage0_col47[7] = pp[7][33];
        stage0_col47[8] = pp[8][31];
        stage0_col47[9] = pp[9][29];
        stage0_col47[10] = pp[10][27];
        stage0_col47[11] = pp[11][25];
        stage0_col47[12] = pp[12][23];
        stage0_col47[13] = pp[13][21];
        stage0_col47[14] = pp[14][19];
        stage0_col47[15] = pp[15][17];
        stage0_col47[16] = pp[16][15];
        stage0_col47[17] = pp[17][13];
        stage0_col47[18] = pp[18][11];
        stage0_col47[19] = pp[19][9];
        stage0_col47[20] = pp[20][7];
        stage0_col47[21] = pp[21][5];
        stage0_col47[22] = pp[22][3];
        stage0_col47[23] = pp[23][1];
        stage0_col48[0] = pp[0][48];
        stage0_col48[1] = pp[1][46];
        stage0_col48[2] = pp[2][44];
        stage0_col48[3] = pp[3][42];
        stage0_col48[4] = pp[4][40];
        stage0_col48[5] = pp[5][38];
        stage0_col48[6] = pp[6][36];
        stage0_col48[7] = pp[7][34];
        stage0_col48[8] = pp[8][32];
        stage0_col48[9] = pp[9][30];
        stage0_col48[10] = pp[10][28];
        stage0_col48[11] = pp[11][26];
        stage0_col48[12] = pp[12][24];
        stage0_col48[13] = pp[13][22];
        stage0_col48[14] = pp[14][20];
        stage0_col48[15] = pp[15][18];
        stage0_col48[16] = pp[16][16];
        stage0_col48[17] = pp[17][14];
        stage0_col48[18] = pp[18][12];
        stage0_col48[19] = pp[19][10];
        stage0_col48[20] = pp[20][8];
        stage0_col48[21] = pp[21][6];
        stage0_col48[22] = pp[22][4];
        stage0_col48[23] = pp[23][2];
        stage0_col48[24] = cpl[24];
        stage0_col48[25] = pp[24][0];
        stage0_col49[0] = pp[0][49];
        stage0_col49[1] = pp[1][47];
        stage0_col49[2] = pp[2][45];
        stage0_col49[3] = pp[3][43];
        stage0_col49[4] = pp[4][41];
        stage0_col49[5] = pp[5][39];
        stage0_col49[6] = pp[6][37];
        stage0_col49[7] = pp[7][35];
        stage0_col49[8] = pp[8][33];
        stage0_col49[9] = pp[9][31];
        stage0_col49[10] = pp[10][29];
        stage0_col49[11] = pp[11][27];
        stage0_col49[12] = pp[12][25];
        stage0_col49[13] = pp[13][23];
        stage0_col49[14] = pp[14][21];
        stage0_col49[15] = pp[15][19];
        stage0_col49[16] = pp[16][17];
        stage0_col49[17] = pp[17][15];
        stage0_col49[18] = pp[18][13];
        stage0_col49[19] = pp[19][11];
        stage0_col49[20] = pp[20][9];
        stage0_col49[21] = pp[21][7];
        stage0_col49[22] = pp[22][5];
        stage0_col49[23] = pp[23][3];
        stage0_col49[24] = pp[24][1];
        stage0_col50[0] = pp[0][50];
        stage0_col50[1] = pp[1][48];
        stage0_col50[2] = pp[2][46];
        stage0_col50[3] = pp[3][44];
        stage0_col50[4] = pp[4][42];
        stage0_col50[5] = pp[5][40];
        stage0_col50[6] = pp[6][38];
        stage0_col50[7] = pp[7][36];
        stage0_col50[8] = pp[8][34];
        stage0_col50[9] = pp[9][32];
        stage0_col50[10] = pp[10][30];
        stage0_col50[11] = pp[11][28];
        stage0_col50[12] = pp[12][26];
        stage0_col50[13] = pp[13][24];
        stage0_col50[14] = pp[14][22];
        stage0_col50[15] = pp[15][20];
        stage0_col50[16] = pp[16][18];
        stage0_col50[17] = pp[17][16];
        stage0_col50[18] = pp[18][14];
        stage0_col50[19] = pp[19][12];
        stage0_col50[20] = pp[20][10];
        stage0_col50[21] = pp[21][8];
        stage0_col50[22] = pp[22][6];
        stage0_col50[23] = pp[23][4];
        stage0_col50[24] = pp[24][2];
        stage0_col50[25] = cpl[25];
        stage0_col50[26] = pp[25][0];
        stage0_col51[0] = pp[0][51];
        stage0_col51[1] = pp[1][49];
        stage0_col51[2] = pp[2][47];
        stage0_col51[3] = pp[3][45];
        stage0_col51[4] = pp[4][43];
        stage0_col51[5] = pp[5][41];
        stage0_col51[6] = pp[6][39];
        stage0_col51[7] = pp[7][37];
        stage0_col51[8] = pp[8][35];
        stage0_col51[9] = pp[9][33];
        stage0_col51[10] = pp[10][31];
        stage0_col51[11] = pp[11][29];
        stage0_col51[12] = pp[12][27];
        stage0_col51[13] = pp[13][25];
        stage0_col51[14] = pp[14][23];
        stage0_col51[15] = pp[15][21];
        stage0_col51[16] = pp[16][19];
        stage0_col51[17] = pp[17][17];
        stage0_col51[18] = pp[18][15];
        stage0_col51[19] = pp[19][13];
        stage0_col51[20] = pp[20][11];
        stage0_col51[21] = pp[21][9];
        stage0_col51[22] = pp[22][7];
        stage0_col51[23] = pp[23][5];
        stage0_col51[24] = pp[24][3];
        stage0_col51[25] = pp[25][1];
        stage0_col52[0] = pp[0][52];
        stage0_col52[1] = pp[1][50];
        stage0_col52[2] = pp[2][48];
        stage0_col52[3] = pp[3][46];
        stage0_col52[4] = pp[4][44];
        stage0_col52[5] = pp[5][42];
        stage0_col52[6] = pp[6][40];
        stage0_col52[7] = pp[7][38];
        stage0_col52[8] = pp[8][36];
        stage0_col52[9] = pp[9][34];
        stage0_col52[10] = pp[10][32];
        stage0_col52[11] = pp[11][30];
        stage0_col52[12] = pp[12][28];
        stage0_col52[13] = pp[13][26];
        stage0_col52[14] = pp[14][24];
        stage0_col52[15] = pp[15][22];
        stage0_col52[16] = pp[16][20];
        stage0_col52[17] = pp[17][18];
        stage0_col52[18] = pp[18][16];
        stage0_col52[19] = pp[19][14];
        stage0_col52[20] = pp[20][12];
        stage0_col52[21] = pp[21][10];
        stage0_col52[22] = pp[22][8];
        stage0_col52[23] = pp[23][6];
        stage0_col52[24] = pp[24][4];
        stage0_col52[25] = pp[25][2];
        stage0_col52[26] = cpl[26];
        stage0_col52[27] = pp[26][0];
        stage0_col53[0] = pp[0][53];
        stage0_col53[1] = pp[1][51];
        stage0_col53[2] = pp[2][49];
        stage0_col53[3] = pp[3][47];
        stage0_col53[4] = pp[4][45];
        stage0_col53[5] = pp[5][43];
        stage0_col53[6] = pp[6][41];
        stage0_col53[7] = pp[7][39];
        stage0_col53[8] = pp[8][37];
        stage0_col53[9] = pp[9][35];
        stage0_col53[10] = pp[10][33];
        stage0_col53[11] = pp[11][31];
        stage0_col53[12] = pp[12][29];
        stage0_col53[13] = pp[13][27];
        stage0_col53[14] = pp[14][25];
        stage0_col53[15] = pp[15][23];
        stage0_col53[16] = pp[16][21];
        stage0_col53[17] = pp[17][19];
        stage0_col53[18] = pp[18][17];
        stage0_col53[19] = pp[19][15];
        stage0_col53[20] = pp[20][13];
        stage0_col53[21] = pp[21][11];
        stage0_col53[22] = pp[22][9];
        stage0_col53[23] = pp[23][7];
        stage0_col53[24] = pp[24][5];
        stage0_col53[25] = pp[25][3];
        stage0_col53[26] = pp[26][1];
        stage0_col54[0] = pp[0][54];
        stage0_col54[1] = pp[1][52];
        stage0_col54[2] = pp[2][50];
        stage0_col54[3] = pp[3][48];
        stage0_col54[4] = pp[4][46];
        stage0_col54[5] = pp[5][44];
        stage0_col54[6] = pp[6][42];
        stage0_col54[7] = pp[7][40];
        stage0_col54[8] = pp[8][38];
        stage0_col54[9] = pp[9][36];
        stage0_col54[10] = pp[10][34];
        stage0_col54[11] = pp[11][32];
        stage0_col54[12] = pp[12][30];
        stage0_col54[13] = pp[13][28];
        stage0_col54[14] = pp[14][26];
        stage0_col54[15] = pp[15][24];
        stage0_col54[16] = pp[16][22];
        stage0_col54[17] = pp[17][20];
        stage0_col54[18] = pp[18][18];
        stage0_col54[19] = pp[19][16];
        stage0_col54[20] = pp[20][14];
        stage0_col54[21] = pp[21][12];
        stage0_col54[22] = pp[22][10];
        stage0_col54[23] = pp[23][8];
        stage0_col54[24] = pp[24][6];
        stage0_col54[25] = pp[25][4];
        stage0_col54[26] = pp[26][2];
        stage0_col54[27] = cpl[27];
        stage0_col54[28] = pp[27][0];
        stage0_col55[0] = pp[0][55];
        stage0_col55[1] = pp[1][53];
        stage0_col55[2] = pp[2][51];
        stage0_col55[3] = pp[3][49];
        stage0_col55[4] = pp[4][47];
        stage0_col55[5] = pp[5][45];
        stage0_col55[6] = pp[6][43];
        stage0_col55[7] = pp[7][41];
        stage0_col55[8] = pp[8][39];
        stage0_col55[9] = pp[9][37];
        stage0_col55[10] = pp[10][35];
        stage0_col55[11] = pp[11][33];
        stage0_col55[12] = pp[12][31];
        stage0_col55[13] = pp[13][29];
        stage0_col55[14] = pp[14][27];
        stage0_col55[15] = pp[15][25];
        stage0_col55[16] = pp[16][23];
        stage0_col55[17] = pp[17][21];
        stage0_col55[18] = pp[18][19];
        stage0_col55[19] = pp[19][17];
        stage0_col55[20] = pp[20][15];
        stage0_col55[21] = pp[21][13];
        stage0_col55[22] = pp[22][11];
        stage0_col55[23] = pp[23][9];
        stage0_col55[24] = pp[24][7];
        stage0_col55[25] = pp[25][5];
        stage0_col55[26] = pp[26][3];
        stage0_col55[27] = pp[27][1];
        stage0_col56[0] = pp[0][56];
        stage0_col56[1] = pp[1][54];
        stage0_col56[2] = pp[2][52];
        stage0_col56[3] = pp[3][50];
        stage0_col56[4] = pp[4][48];
        stage0_col56[5] = pp[5][46];
        stage0_col56[6] = pp[6][44];
        stage0_col56[7] = pp[7][42];
        stage0_col56[8] = pp[8][40];
        stage0_col56[9] = pp[9][38];
        stage0_col56[10] = pp[10][36];
        stage0_col56[11] = pp[11][34];
        stage0_col56[12] = pp[12][32];
        stage0_col56[13] = pp[13][30];
        stage0_col56[14] = pp[14][28];
        stage0_col56[15] = pp[15][26];
        stage0_col56[16] = pp[16][24];
        stage0_col56[17] = pp[17][22];
        stage0_col56[18] = pp[18][20];
        stage0_col56[19] = pp[19][18];
        stage0_col56[20] = pp[20][16];
        stage0_col56[21] = pp[21][14];
        stage0_col56[22] = pp[22][12];
        stage0_col56[23] = pp[23][10];
        stage0_col56[24] = pp[24][8];
        stage0_col56[25] = pp[25][6];
        stage0_col56[26] = pp[26][4];
        stage0_col56[27] = pp[27][2];
        stage0_col56[28] = cpl[28];
        stage0_col56[29] = pp[28][0];
        stage0_col57[0] = pp[0][57];
        stage0_col57[1] = pp[1][55];
        stage0_col57[2] = pp[2][53];
        stage0_col57[3] = pp[3][51];
        stage0_col57[4] = pp[4][49];
        stage0_col57[5] = pp[5][47];
        stage0_col57[6] = pp[6][45];
        stage0_col57[7] = pp[7][43];
        stage0_col57[8] = pp[8][41];
        stage0_col57[9] = pp[9][39];
        stage0_col57[10] = pp[10][37];
        stage0_col57[11] = pp[11][35];
        stage0_col57[12] = pp[12][33];
        stage0_col57[13] = pp[13][31];
        stage0_col57[14] = pp[14][29];
        stage0_col57[15] = pp[15][27];
        stage0_col57[16] = pp[16][25];
        stage0_col57[17] = pp[17][23];
        stage0_col57[18] = pp[18][21];
        stage0_col57[19] = pp[19][19];
        stage0_col57[20] = pp[20][17];
        stage0_col57[21] = pp[21][15];
        stage0_col57[22] = pp[22][13];
        stage0_col57[23] = pp[23][11];
        stage0_col57[24] = pp[24][9];
        stage0_col57[25] = pp[25][7];
        stage0_col57[26] = pp[26][5];
        stage0_col57[27] = pp[27][3];
        stage0_col57[28] = pp[28][1];
        stage0_col58[0] = pp[0][58];
        stage0_col58[1] = pp[1][56];
        stage0_col58[2] = pp[2][54];
        stage0_col58[3] = pp[3][52];
        stage0_col58[4] = pp[4][50];
        stage0_col58[5] = pp[5][48];
        stage0_col58[6] = pp[6][46];
        stage0_col58[7] = pp[7][44];
        stage0_col58[8] = pp[8][42];
        stage0_col58[9] = pp[9][40];
        stage0_col58[10] = pp[10][38];
        stage0_col58[11] = pp[11][36];
        stage0_col58[12] = pp[12][34];
        stage0_col58[13] = pp[13][32];
        stage0_col58[14] = pp[14][30];
        stage0_col58[15] = pp[15][28];
        stage0_col58[16] = pp[16][26];
        stage0_col58[17] = pp[17][24];
        stage0_col58[18] = pp[18][22];
        stage0_col58[19] = pp[19][20];
        stage0_col58[20] = pp[20][18];
        stage0_col58[21] = pp[21][16];
        stage0_col58[22] = pp[22][14];
        stage0_col58[23] = pp[23][12];
        stage0_col58[24] = pp[24][10];
        stage0_col58[25] = pp[25][8];
        stage0_col58[26] = pp[26][6];
        stage0_col58[27] = pp[27][4];
        stage0_col58[28] = pp[28][2];
        stage0_col58[29] = cpl[29];
        stage0_col58[30] = pp[29][0];
        stage0_col59[0] = pp[0][59];
        stage0_col59[1] = pp[1][57];
        stage0_col59[2] = pp[2][55];
        stage0_col59[3] = pp[3][53];
        stage0_col59[4] = pp[4][51];
        stage0_col59[5] = pp[5][49];
        stage0_col59[6] = pp[6][47];
        stage0_col59[7] = pp[7][45];
        stage0_col59[8] = pp[8][43];
        stage0_col59[9] = pp[9][41];
        stage0_col59[10] = pp[10][39];
        stage0_col59[11] = pp[11][37];
        stage0_col59[12] = pp[12][35];
        stage0_col59[13] = pp[13][33];
        stage0_col59[14] = pp[14][31];
        stage0_col59[15] = pp[15][29];
        stage0_col59[16] = pp[16][27];
        stage0_col59[17] = pp[17][25];
        stage0_col59[18] = pp[18][23];
        stage0_col59[19] = pp[19][21];
        stage0_col59[20] = pp[20][19];
        stage0_col59[21] = pp[21][17];
        stage0_col59[22] = pp[22][15];
        stage0_col59[23] = pp[23][13];
        stage0_col59[24] = pp[24][11];
        stage0_col59[25] = pp[25][9];
        stage0_col59[26] = pp[26][7];
        stage0_col59[27] = pp[27][5];
        stage0_col59[28] = pp[28][3];
        stage0_col59[29] = pp[29][1];
        stage0_col60[0] = pp[0][60];
        stage0_col60[1] = pp[1][58];
        stage0_col60[2] = pp[2][56];
        stage0_col60[3] = pp[3][54];
        stage0_col60[4] = pp[4][52];
        stage0_col60[5] = pp[5][50];
        stage0_col60[6] = pp[6][48];
        stage0_col60[7] = pp[7][46];
        stage0_col60[8] = pp[8][44];
        stage0_col60[9] = pp[9][42];
        stage0_col60[10] = pp[10][40];
        stage0_col60[11] = pp[11][38];
        stage0_col60[12] = pp[12][36];
        stage0_col60[13] = pp[13][34];
        stage0_col60[14] = pp[14][32];
        stage0_col60[15] = pp[15][30];
        stage0_col60[16] = pp[16][28];
        stage0_col60[17] = pp[17][26];
        stage0_col60[18] = pp[18][24];
        stage0_col60[19] = pp[19][22];
        stage0_col60[20] = pp[20][20];
        stage0_col60[21] = pp[21][18];
        stage0_col60[22] = pp[22][16];
        stage0_col60[23] = pp[23][14];
        stage0_col60[24] = pp[24][12];
        stage0_col60[25] = pp[25][10];
        stage0_col60[26] = pp[26][8];
        stage0_col60[27] = pp[27][6];
        stage0_col60[28] = pp[28][4];
        stage0_col60[29] = pp[29][2];
        stage0_col60[30] = cpl[30];
        stage0_col60[31] = pp[30][0];
        stage0_col61[0] = pp[0][61];
        stage0_col61[1] = pp[1][59];
        stage0_col61[2] = pp[2][57];
        stage0_col61[3] = pp[3][55];
        stage0_col61[4] = pp[4][53];
        stage0_col61[5] = pp[5][51];
        stage0_col61[6] = pp[6][49];
        stage0_col61[7] = pp[7][47];
        stage0_col61[8] = pp[8][45];
        stage0_col61[9] = pp[9][43];
        stage0_col61[10] = pp[10][41];
        stage0_col61[11] = pp[11][39];
        stage0_col61[12] = pp[12][37];
        stage0_col61[13] = pp[13][35];
        stage0_col61[14] = pp[14][33];
        stage0_col61[15] = pp[15][31];
        stage0_col61[16] = pp[16][29];
        stage0_col61[17] = pp[17][27];
        stage0_col61[18] = pp[18][25];
        stage0_col61[19] = pp[19][23];
        stage0_col61[20] = pp[20][21];
        stage0_col61[21] = pp[21][19];
        stage0_col61[22] = pp[22][17];
        stage0_col61[23] = pp[23][15];
        stage0_col61[24] = pp[24][13];
        stage0_col61[25] = pp[25][11];
        stage0_col61[26] = pp[26][9];
        stage0_col61[27] = pp[27][7];
        stage0_col61[28] = pp[28][5];
        stage0_col61[29] = pp[29][3];
        stage0_col61[30] = pp[30][1];
        stage0_col62[0] = pp[0][62];
        stage0_col62[1] = pp[1][60];
        stage0_col62[2] = pp[2][58];
        stage0_col62[3] = pp[3][56];
        stage0_col62[4] = pp[4][54];
        stage0_col62[5] = pp[5][52];
        stage0_col62[6] = pp[6][50];
        stage0_col62[7] = pp[7][48];
        stage0_col62[8] = pp[8][46];
        stage0_col62[9] = pp[9][44];
        stage0_col62[10] = pp[10][42];
        stage0_col62[11] = pp[11][40];
        stage0_col62[12] = pp[12][38];
        stage0_col62[13] = pp[13][36];
        stage0_col62[14] = pp[14][34];
        stage0_col62[15] = pp[15][32];
        stage0_col62[16] = pp[16][30];
        stage0_col62[17] = pp[17][28];
        stage0_col62[18] = pp[18][26];
        stage0_col62[19] = pp[19][24];
        stage0_col62[20] = pp[20][22];
        stage0_col62[21] = pp[21][20];
        stage0_col62[22] = pp[22][18];
        stage0_col62[23] = pp[23][16];
        stage0_col62[24] = pp[24][14];
        stage0_col62[25] = pp[25][12];
        stage0_col62[26] = pp[26][10];
        stage0_col62[27] = pp[27][8];
        stage0_col62[28] = pp[28][6];
        stage0_col62[29] = pp[29][4];
        stage0_col62[30] = pp[30][2];
        stage0_col62[31] = cpl[31];
        stage0_col62[32] = pp[31][0];
        stage0_col63[0] = pp[0][63];
        stage0_col63[1] = pp[1][61];
        stage0_col63[2] = pp[2][59];
        stage0_col63[3] = pp[3][57];
        stage0_col63[4] = pp[4][55];
        stage0_col63[5] = pp[5][53];
        stage0_col63[6] = pp[6][51];
        stage0_col63[7] = pp[7][49];
        stage0_col63[8] = pp[8][47];
        stage0_col63[9] = pp[9][45];
        stage0_col63[10] = pp[10][43];
        stage0_col63[11] = pp[11][41];
        stage0_col63[12] = pp[12][39];
        stage0_col63[13] = pp[13][37];
        stage0_col63[14] = pp[14][35];
        stage0_col63[15] = pp[15][33];
        stage0_col63[16] = pp[16][31];
        stage0_col63[17] = pp[17][29];
        stage0_col63[18] = pp[18][27];
        stage0_col63[19] = pp[19][25];
        stage0_col63[20] = pp[20][23];
        stage0_col63[21] = pp[21][21];
        stage0_col63[22] = pp[22][19];
        stage0_col63[23] = pp[23][17];
        stage0_col63[24] = pp[24][15];
        stage0_col63[25] = pp[25][13];
        stage0_col63[26] = pp[26][11];
        stage0_col63[27] = pp[27][9];
        stage0_col63[28] = pp[28][7];
        stage0_col63[29] = pp[29][5];
        stage0_col63[30] = pp[30][3];
        stage0_col63[31] = pp[31][1];
        stage0_col64[0] = ~pp[0][64];
        stage0_col64[1] = 1'b1;
        stage0_col64[2] = pp[1][62];
        stage0_col64[3] = pp[2][60];
        stage0_col64[4] = pp[3][58];
        stage0_col64[5] = pp[4][56];
        stage0_col64[6] = pp[5][54];
        stage0_col64[7] = pp[6][52];
        stage0_col64[8] = pp[7][50];
        stage0_col64[9] = pp[8][48];
        stage0_col64[10] = pp[9][46];
        stage0_col64[11] = pp[10][44];
        stage0_col64[12] = pp[11][42];
        stage0_col64[13] = pp[12][40];
        stage0_col64[14] = pp[13][38];
        stage0_col64[15] = pp[14][36];
        stage0_col64[16] = pp[15][34];
        stage0_col64[17] = pp[16][32];
        stage0_col64[18] = pp[17][30];
        stage0_col64[19] = pp[18][28];
        stage0_col64[20] = pp[19][26];
        stage0_col64[21] = pp[20][24];
        stage0_col64[22] = pp[21][22];
        stage0_col64[23] = pp[22][20];
        stage0_col64[24] = pp[23][18];
        stage0_col64[25] = pp[24][16];
        stage0_col64[26] = pp[25][14];
        stage0_col64[27] = pp[26][12];
        stage0_col64[28] = pp[27][10];
        stage0_col64[29] = pp[28][8];
        stage0_col64[30] = pp[29][6];
        stage0_col64[31] = pp[30][4];
        stage0_col64[32] = pp[31][2];
        stage0_col65[0] = 1'b1;
        stage0_col65[1] = pp[1][63];
        stage0_col65[2] = pp[2][61];
        stage0_col65[3] = pp[3][59];
        stage0_col65[4] = pp[4][57];
        stage0_col65[5] = pp[5][55];
        stage0_col65[6] = pp[6][53];
        stage0_col65[7] = pp[7][51];
        stage0_col65[8] = pp[8][49];
        stage0_col65[9] = pp[9][47];
        stage0_col65[10] = pp[10][45];
        stage0_col65[11] = pp[11][43];
        stage0_col65[12] = pp[12][41];
        stage0_col65[13] = pp[13][39];
        stage0_col65[14] = pp[14][37];
        stage0_col65[15] = pp[15][35];
        stage0_col65[16] = pp[16][33];
        stage0_col65[17] = pp[17][31];
        stage0_col65[18] = pp[18][29];
        stage0_col65[19] = pp[19][27];
        stage0_col65[20] = pp[20][25];
        stage0_col65[21] = pp[21][23];
        stage0_col65[22] = pp[22][21];
        stage0_col65[23] = pp[23][19];
        stage0_col65[24] = pp[24][17];
        stage0_col65[25] = pp[25][15];
        stage0_col65[26] = pp[26][13];
        stage0_col65[27] = pp[27][11];
        stage0_col65[28] = pp[28][9];
        stage0_col65[29] = pp[29][7];
        stage0_col65[30] = pp[30][5];
        stage0_col65[31] = pp[31][3];
        stage0_col66[0] = 1'b1;
        stage0_col66[1] = ~pp[1][64];
        stage0_col66[2] = 1'b1;
        stage0_col66[3] = pp[2][62];
        stage0_col66[4] = pp[3][60];
        stage0_col66[5] = pp[4][58];
        stage0_col66[6] = pp[5][56];
        stage0_col66[7] = pp[6][54];
        stage0_col66[8] = pp[7][52];
        stage0_col66[9] = pp[8][50];
        stage0_col66[10] = pp[9][48];
        stage0_col66[11] = pp[10][46];
        stage0_col66[12] = pp[11][44];
        stage0_col66[13] = pp[12][42];
        stage0_col66[14] = pp[13][40];
        stage0_col66[15] = pp[14][38];
        stage0_col66[16] = pp[15][36];
        stage0_col66[17] = pp[16][34];
        stage0_col66[18] = pp[17][32];
        stage0_col66[19] = pp[18][30];
        stage0_col66[20] = pp[19][28];
        stage0_col66[21] = pp[20][26];
        stage0_col66[22] = pp[21][24];
        stage0_col66[23] = pp[22][22];
        stage0_col66[24] = pp[23][20];
        stage0_col66[25] = pp[24][18];
        stage0_col66[26] = pp[25][16];
        stage0_col66[27] = pp[26][14];
        stage0_col66[28] = pp[27][12];
        stage0_col66[29] = pp[28][10];
        stage0_col66[30] = pp[29][8];
        stage0_col66[31] = pp[30][6];
        stage0_col66[32] = pp[31][4];
        stage0_col67[0] = 1'b1;
        stage0_col67[1] = 1'b1;
        stage0_col67[2] = pp[2][63];
        stage0_col67[3] = pp[3][61];
        stage0_col67[4] = pp[4][59];
        stage0_col67[5] = pp[5][57];
        stage0_col67[6] = pp[6][55];
        stage0_col67[7] = pp[7][53];
        stage0_col67[8] = pp[8][51];
        stage0_col67[9] = pp[9][49];
        stage0_col67[10] = pp[10][47];
        stage0_col67[11] = pp[11][45];
        stage0_col67[12] = pp[12][43];
        stage0_col67[13] = pp[13][41];
        stage0_col67[14] = pp[14][39];
        stage0_col67[15] = pp[15][37];
        stage0_col67[16] = pp[16][35];
        stage0_col67[17] = pp[17][33];
        stage0_col67[18] = pp[18][31];
        stage0_col67[19] = pp[19][29];
        stage0_col67[20] = pp[20][27];
        stage0_col67[21] = pp[21][25];
        stage0_col67[22] = pp[22][23];
        stage0_col67[23] = pp[23][21];
        stage0_col67[24] = pp[24][19];
        stage0_col67[25] = pp[25][17];
        stage0_col67[26] = pp[26][15];
        stage0_col67[27] = pp[27][13];
        stage0_col67[28] = pp[28][11];
        stage0_col67[29] = pp[29][9];
        stage0_col67[30] = pp[30][7];
        stage0_col67[31] = pp[31][5];
        stage0_col68[0] = 1'b1;
        stage0_col68[1] = 1'b1;
        stage0_col68[2] = ~pp[2][64];
        stage0_col68[3] = 1'b1;
        stage0_col68[4] = pp[3][62];
        stage0_col68[5] = pp[4][60];
        stage0_col68[6] = pp[5][58];
        stage0_col68[7] = pp[6][56];
        stage0_col68[8] = pp[7][54];
        stage0_col68[9] = pp[8][52];
        stage0_col68[10] = pp[9][50];
        stage0_col68[11] = pp[10][48];
        stage0_col68[12] = pp[11][46];
        stage0_col68[13] = pp[12][44];
        stage0_col68[14] = pp[13][42];
        stage0_col68[15] = pp[14][40];
        stage0_col68[16] = pp[15][38];
        stage0_col68[17] = pp[16][36];
        stage0_col68[18] = pp[17][34];
        stage0_col68[19] = pp[18][32];
        stage0_col68[20] = pp[19][30];
        stage0_col68[21] = pp[20][28];
        stage0_col68[22] = pp[21][26];
        stage0_col68[23] = pp[22][24];
        stage0_col68[24] = pp[23][22];
        stage0_col68[25] = pp[24][20];
        stage0_col68[26] = pp[25][18];
        stage0_col68[27] = pp[26][16];
        stage0_col68[28] = pp[27][14];
        stage0_col68[29] = pp[28][12];
        stage0_col68[30] = pp[29][10];
        stage0_col68[31] = pp[30][8];
        stage0_col68[32] = pp[31][6];
        stage0_col69[0] = 1'b1;
        stage0_col69[1] = 1'b1;
        stage0_col69[2] = 1'b1;
        stage0_col69[3] = pp[3][63];
        stage0_col69[4] = pp[4][61];
        stage0_col69[5] = pp[5][59];
        stage0_col69[6] = pp[6][57];
        stage0_col69[7] = pp[7][55];
        stage0_col69[8] = pp[8][53];
        stage0_col69[9] = pp[9][51];
        stage0_col69[10] = pp[10][49];
        stage0_col69[11] = pp[11][47];
        stage0_col69[12] = pp[12][45];
        stage0_col69[13] = pp[13][43];
        stage0_col69[14] = pp[14][41];
        stage0_col69[15] = pp[15][39];
        stage0_col69[16] = pp[16][37];
        stage0_col69[17] = pp[17][35];
        stage0_col69[18] = pp[18][33];
        stage0_col69[19] = pp[19][31];
        stage0_col69[20] = pp[20][29];
        stage0_col69[21] = pp[21][27];
        stage0_col69[22] = pp[22][25];
        stage0_col69[23] = pp[23][23];
        stage0_col69[24] = pp[24][21];
        stage0_col69[25] = pp[25][19];
        stage0_col69[26] = pp[26][17];
        stage0_col69[27] = pp[27][15];
        stage0_col69[28] = pp[28][13];
        stage0_col69[29] = pp[29][11];
        stage0_col69[30] = pp[30][9];
        stage0_col69[31] = pp[31][7];
        stage0_col70[0] = 1'b1;
        stage0_col70[1] = 1'b1;
        stage0_col70[2] = 1'b1;
        stage0_col70[3] = ~pp[3][64];
        stage0_col70[4] = 1'b1;
        stage0_col70[5] = pp[4][62];
        stage0_col70[6] = pp[5][60];
        stage0_col70[7] = pp[6][58];
        stage0_col70[8] = pp[7][56];
        stage0_col70[9] = pp[8][54];
        stage0_col70[10] = pp[9][52];
        stage0_col70[11] = pp[10][50];
        stage0_col70[12] = pp[11][48];
        stage0_col70[13] = pp[12][46];
        stage0_col70[14] = pp[13][44];
        stage0_col70[15] = pp[14][42];
        stage0_col70[16] = pp[15][40];
        stage0_col70[17] = pp[16][38];
        stage0_col70[18] = pp[17][36];
        stage0_col70[19] = pp[18][34];
        stage0_col70[20] = pp[19][32];
        stage0_col70[21] = pp[20][30];
        stage0_col70[22] = pp[21][28];
        stage0_col70[23] = pp[22][26];
        stage0_col70[24] = pp[23][24];
        stage0_col70[25] = pp[24][22];
        stage0_col70[26] = pp[25][20];
        stage0_col70[27] = pp[26][18];
        stage0_col70[28] = pp[27][16];
        stage0_col70[29] = pp[28][14];
        stage0_col70[30] = pp[29][12];
        stage0_col70[31] = pp[30][10];
        stage0_col70[32] = pp[31][8];
        stage0_col71[0] = 1'b1;
        stage0_col71[1] = 1'b1;
        stage0_col71[2] = 1'b1;
        stage0_col71[3] = 1'b1;
        stage0_col71[4] = pp[4][63];
        stage0_col71[5] = pp[5][61];
        stage0_col71[6] = pp[6][59];
        stage0_col71[7] = pp[7][57];
        stage0_col71[8] = pp[8][55];
        stage0_col71[9] = pp[9][53];
        stage0_col71[10] = pp[10][51];
        stage0_col71[11] = pp[11][49];
        stage0_col71[12] = pp[12][47];
        stage0_col71[13] = pp[13][45];
        stage0_col71[14] = pp[14][43];
        stage0_col71[15] = pp[15][41];
        stage0_col71[16] = pp[16][39];
        stage0_col71[17] = pp[17][37];
        stage0_col71[18] = pp[18][35];
        stage0_col71[19] = pp[19][33];
        stage0_col71[20] = pp[20][31];
        stage0_col71[21] = pp[21][29];
        stage0_col71[22] = pp[22][27];
        stage0_col71[23] = pp[23][25];
        stage0_col71[24] = pp[24][23];
        stage0_col71[25] = pp[25][21];
        stage0_col71[26] = pp[26][19];
        stage0_col71[27] = pp[27][17];
        stage0_col71[28] = pp[28][15];
        stage0_col71[29] = pp[29][13];
        stage0_col71[30] = pp[30][11];
        stage0_col71[31] = pp[31][9];
        stage0_col72[0] = 1'b1;
        stage0_col72[1] = 1'b1;
        stage0_col72[2] = 1'b1;
        stage0_col72[3] = 1'b1;
        stage0_col72[4] = ~pp[4][64];
        stage0_col72[5] = 1'b1;
        stage0_col72[6] = pp[5][62];
        stage0_col72[7] = pp[6][60];
        stage0_col72[8] = pp[7][58];
        stage0_col72[9] = pp[8][56];
        stage0_col72[10] = pp[9][54];
        stage0_col72[11] = pp[10][52];
        stage0_col72[12] = pp[11][50];
        stage0_col72[13] = pp[12][48];
        stage0_col72[14] = pp[13][46];
        stage0_col72[15] = pp[14][44];
        stage0_col72[16] = pp[15][42];
        stage0_col72[17] = pp[16][40];
        stage0_col72[18] = pp[17][38];
        stage0_col72[19] = pp[18][36];
        stage0_col72[20] = pp[19][34];
        stage0_col72[21] = pp[20][32];
        stage0_col72[22] = pp[21][30];
        stage0_col72[23] = pp[22][28];
        stage0_col72[24] = pp[23][26];
        stage0_col72[25] = pp[24][24];
        stage0_col72[26] = pp[25][22];
        stage0_col72[27] = pp[26][20];
        stage0_col72[28] = pp[27][18];
        stage0_col72[29] = pp[28][16];
        stage0_col72[30] = pp[29][14];
        stage0_col72[31] = pp[30][12];
        stage0_col72[32] = pp[31][10];
        stage0_col73[0] = 1'b1;
        stage0_col73[1] = 1'b1;
        stage0_col73[2] = 1'b1;
        stage0_col73[3] = 1'b1;
        stage0_col73[4] = 1'b1;
        stage0_col73[5] = pp[5][63];
        stage0_col73[6] = pp[6][61];
        stage0_col73[7] = pp[7][59];
        stage0_col73[8] = pp[8][57];
        stage0_col73[9] = pp[9][55];
        stage0_col73[10] = pp[10][53];
        stage0_col73[11] = pp[11][51];
        stage0_col73[12] = pp[12][49];
        stage0_col73[13] = pp[13][47];
        stage0_col73[14] = pp[14][45];
        stage0_col73[15] = pp[15][43];
        stage0_col73[16] = pp[16][41];
        stage0_col73[17] = pp[17][39];
        stage0_col73[18] = pp[18][37];
        stage0_col73[19] = pp[19][35];
        stage0_col73[20] = pp[20][33];
        stage0_col73[21] = pp[21][31];
        stage0_col73[22] = pp[22][29];
        stage0_col73[23] = pp[23][27];
        stage0_col73[24] = pp[24][25];
        stage0_col73[25] = pp[25][23];
        stage0_col73[26] = pp[26][21];
        stage0_col73[27] = pp[27][19];
        stage0_col73[28] = pp[28][17];
        stage0_col73[29] = pp[29][15];
        stage0_col73[30] = pp[30][13];
        stage0_col73[31] = pp[31][11];
        stage0_col74[0] = 1'b1;
        stage0_col74[1] = 1'b1;
        stage0_col74[2] = 1'b1;
        stage0_col74[3] = 1'b1;
        stage0_col74[4] = 1'b1;
        stage0_col74[5] = ~pp[5][64];
        stage0_col74[6] = 1'b1;
        stage0_col74[7] = pp[6][62];
        stage0_col74[8] = pp[7][60];
        stage0_col74[9] = pp[8][58];
        stage0_col74[10] = pp[9][56];
        stage0_col74[11] = pp[10][54];
        stage0_col74[12] = pp[11][52];
        stage0_col74[13] = pp[12][50];
        stage0_col74[14] = pp[13][48];
        stage0_col74[15] = pp[14][46];
        stage0_col74[16] = pp[15][44];
        stage0_col74[17] = pp[16][42];
        stage0_col74[18] = pp[17][40];
        stage0_col74[19] = pp[18][38];
        stage0_col74[20] = pp[19][36];
        stage0_col74[21] = pp[20][34];
        stage0_col74[22] = pp[21][32];
        stage0_col74[23] = pp[22][30];
        stage0_col74[24] = pp[23][28];
        stage0_col74[25] = pp[24][26];
        stage0_col74[26] = pp[25][24];
        stage0_col74[27] = pp[26][22];
        stage0_col74[28] = pp[27][20];
        stage0_col74[29] = pp[28][18];
        stage0_col74[30] = pp[29][16];
        stage0_col74[31] = pp[30][14];
        stage0_col74[32] = pp[31][12];
        stage0_col75[0] = 1'b1;
        stage0_col75[1] = 1'b1;
        stage0_col75[2] = 1'b1;
        stage0_col75[3] = 1'b1;
        stage0_col75[4] = 1'b1;
        stage0_col75[5] = 1'b1;
        stage0_col75[6] = pp[6][63];
        stage0_col75[7] = pp[7][61];
        stage0_col75[8] = pp[8][59];
        stage0_col75[9] = pp[9][57];
        stage0_col75[10] = pp[10][55];
        stage0_col75[11] = pp[11][53];
        stage0_col75[12] = pp[12][51];
        stage0_col75[13] = pp[13][49];
        stage0_col75[14] = pp[14][47];
        stage0_col75[15] = pp[15][45];
        stage0_col75[16] = pp[16][43];
        stage0_col75[17] = pp[17][41];
        stage0_col75[18] = pp[18][39];
        stage0_col75[19] = pp[19][37];
        stage0_col75[20] = pp[20][35];
        stage0_col75[21] = pp[21][33];
        stage0_col75[22] = pp[22][31];
        stage0_col75[23] = pp[23][29];
        stage0_col75[24] = pp[24][27];
        stage0_col75[25] = pp[25][25];
        stage0_col75[26] = pp[26][23];
        stage0_col75[27] = pp[27][21];
        stage0_col75[28] = pp[28][19];
        stage0_col75[29] = pp[29][17];
        stage0_col75[30] = pp[30][15];
        stage0_col75[31] = pp[31][13];
        stage0_col76[0] = 1'b1;
        stage0_col76[1] = 1'b1;
        stage0_col76[2] = 1'b1;
        stage0_col76[3] = 1'b1;
        stage0_col76[4] = 1'b1;
        stage0_col76[5] = 1'b1;
        stage0_col76[6] = ~pp[6][64];
        stage0_col76[7] = 1'b1;
        stage0_col76[8] = pp[7][62];
        stage0_col76[9] = pp[8][60];
        stage0_col76[10] = pp[9][58];
        stage0_col76[11] = pp[10][56];
        stage0_col76[12] = pp[11][54];
        stage0_col76[13] = pp[12][52];
        stage0_col76[14] = pp[13][50];
        stage0_col76[15] = pp[14][48];
        stage0_col76[16] = pp[15][46];
        stage0_col76[17] = pp[16][44];
        stage0_col76[18] = pp[17][42];
        stage0_col76[19] = pp[18][40];
        stage0_col76[20] = pp[19][38];
        stage0_col76[21] = pp[20][36];
        stage0_col76[22] = pp[21][34];
        stage0_col76[23] = pp[22][32];
        stage0_col76[24] = pp[23][30];
        stage0_col76[25] = pp[24][28];
        stage0_col76[26] = pp[25][26];
        stage0_col76[27] = pp[26][24];
        stage0_col76[28] = pp[27][22];
        stage0_col76[29] = pp[28][20];
        stage0_col76[30] = pp[29][18];
        stage0_col76[31] = pp[30][16];
        stage0_col76[32] = pp[31][14];
        stage0_col77[0] = 1'b1;
        stage0_col77[1] = 1'b1;
        stage0_col77[2] = 1'b1;
        stage0_col77[3] = 1'b1;
        stage0_col77[4] = 1'b1;
        stage0_col77[5] = 1'b1;
        stage0_col77[6] = 1'b1;
        stage0_col77[7] = pp[7][63];
        stage0_col77[8] = pp[8][61];
        stage0_col77[9] = pp[9][59];
        stage0_col77[10] = pp[10][57];
        stage0_col77[11] = pp[11][55];
        stage0_col77[12] = pp[12][53];
        stage0_col77[13] = pp[13][51];
        stage0_col77[14] = pp[14][49];
        stage0_col77[15] = pp[15][47];
        stage0_col77[16] = pp[16][45];
        stage0_col77[17] = pp[17][43];
        stage0_col77[18] = pp[18][41];
        stage0_col77[19] = pp[19][39];
        stage0_col77[20] = pp[20][37];
        stage0_col77[21] = pp[21][35];
        stage0_col77[22] = pp[22][33];
        stage0_col77[23] = pp[23][31];
        stage0_col77[24] = pp[24][29];
        stage0_col77[25] = pp[25][27];
        stage0_col77[26] = pp[26][25];
        stage0_col77[27] = pp[27][23];
        stage0_col77[28] = pp[28][21];
        stage0_col77[29] = pp[29][19];
        stage0_col77[30] = pp[30][17];
        stage0_col77[31] = pp[31][15];
        stage0_col78[0] = 1'b1;
        stage0_col78[1] = 1'b1;
        stage0_col78[2] = 1'b1;
        stage0_col78[3] = 1'b1;
        stage0_col78[4] = 1'b1;
        stage0_col78[5] = 1'b1;
        stage0_col78[6] = 1'b1;
        stage0_col78[7] = ~pp[7][64];
        stage0_col78[8] = 1'b1;
        stage0_col78[9] = pp[8][62];
        stage0_col78[10] = pp[9][60];
        stage0_col78[11] = pp[10][58];
        stage0_col78[12] = pp[11][56];
        stage0_col78[13] = pp[12][54];
        stage0_col78[14] = pp[13][52];
        stage0_col78[15] = pp[14][50];
        stage0_col78[16] = pp[15][48];
        stage0_col78[17] = pp[16][46];
        stage0_col78[18] = pp[17][44];
        stage0_col78[19] = pp[18][42];
        stage0_col78[20] = pp[19][40];
        stage0_col78[21] = pp[20][38];
        stage0_col78[22] = pp[21][36];
        stage0_col78[23] = pp[22][34];
        stage0_col78[24] = pp[23][32];
        stage0_col78[25] = pp[24][30];
        stage0_col78[26] = pp[25][28];
        stage0_col78[27] = pp[26][26];
        stage0_col78[28] = pp[27][24];
        stage0_col78[29] = pp[28][22];
        stage0_col78[30] = pp[29][20];
        stage0_col78[31] = pp[30][18];
        stage0_col78[32] = pp[31][16];
        stage0_col79[0] = 1'b1;
        stage0_col79[1] = 1'b1;
        stage0_col79[2] = 1'b1;
        stage0_col79[3] = 1'b1;
        stage0_col79[4] = 1'b1;
        stage0_col79[5] = 1'b1;
        stage0_col79[6] = 1'b1;
        stage0_col79[7] = 1'b1;
        stage0_col79[8] = pp[8][63];
        stage0_col79[9] = pp[9][61];
        stage0_col79[10] = pp[10][59];
        stage0_col79[11] = pp[11][57];
        stage0_col79[12] = pp[12][55];
        stage0_col79[13] = pp[13][53];
        stage0_col79[14] = pp[14][51];
        stage0_col79[15] = pp[15][49];
        stage0_col79[16] = pp[16][47];
        stage0_col79[17] = pp[17][45];
        stage0_col79[18] = pp[18][43];
        stage0_col79[19] = pp[19][41];
        stage0_col79[20] = pp[20][39];
        stage0_col79[21] = pp[21][37];
        stage0_col79[22] = pp[22][35];
        stage0_col79[23] = pp[23][33];
        stage0_col79[24] = pp[24][31];
        stage0_col79[25] = pp[25][29];
        stage0_col79[26] = pp[26][27];
        stage0_col79[27] = pp[27][25];
        stage0_col79[28] = pp[28][23];
        stage0_col79[29] = pp[29][21];
        stage0_col79[30] = pp[30][19];
        stage0_col79[31] = pp[31][17];
        stage0_col80[0] = 1'b1;
        stage0_col80[1] = 1'b1;
        stage0_col80[2] = 1'b1;
        stage0_col80[3] = 1'b1;
        stage0_col80[4] = 1'b1;
        stage0_col80[5] = 1'b1;
        stage0_col80[6] = 1'b1;
        stage0_col80[7] = 1'b1;
        stage0_col80[8] = ~pp[8][64];
        stage0_col80[9] = 1'b1;
        stage0_col80[10] = pp[9][62];
        stage0_col80[11] = pp[10][60];
        stage0_col80[12] = pp[11][58];
        stage0_col80[13] = pp[12][56];
        stage0_col80[14] = pp[13][54];
        stage0_col80[15] = pp[14][52];
        stage0_col80[16] = pp[15][50];
        stage0_col80[17] = pp[16][48];
        stage0_col80[18] = pp[17][46];
        stage0_col80[19] = pp[18][44];
        stage0_col80[20] = pp[19][42];
        stage0_col80[21] = pp[20][40];
        stage0_col80[22] = pp[21][38];
        stage0_col80[23] = pp[22][36];
        stage0_col80[24] = pp[23][34];
        stage0_col80[25] = pp[24][32];
        stage0_col80[26] = pp[25][30];
        stage0_col80[27] = pp[26][28];
        stage0_col80[28] = pp[27][26];
        stage0_col80[29] = pp[28][24];
        stage0_col80[30] = pp[29][22];
        stage0_col80[31] = pp[30][20];
        stage0_col80[32] = pp[31][18];
        stage0_col81[0] = 1'b1;
        stage0_col81[1] = 1'b1;
        stage0_col81[2] = 1'b1;
        stage0_col81[3] = 1'b1;
        stage0_col81[4] = 1'b1;
        stage0_col81[5] = 1'b1;
        stage0_col81[6] = 1'b1;
        stage0_col81[7] = 1'b1;
        stage0_col81[8] = 1'b1;
        stage0_col81[9] = pp[9][63];
        stage0_col81[10] = pp[10][61];
        stage0_col81[11] = pp[11][59];
        stage0_col81[12] = pp[12][57];
        stage0_col81[13] = pp[13][55];
        stage0_col81[14] = pp[14][53];
        stage0_col81[15] = pp[15][51];
        stage0_col81[16] = pp[16][49];
        stage0_col81[17] = pp[17][47];
        stage0_col81[18] = pp[18][45];
        stage0_col81[19] = pp[19][43];
        stage0_col81[20] = pp[20][41];
        stage0_col81[21] = pp[21][39];
        stage0_col81[22] = pp[22][37];
        stage0_col81[23] = pp[23][35];
        stage0_col81[24] = pp[24][33];
        stage0_col81[25] = pp[25][31];
        stage0_col81[26] = pp[26][29];
        stage0_col81[27] = pp[27][27];
        stage0_col81[28] = pp[28][25];
        stage0_col81[29] = pp[29][23];
        stage0_col81[30] = pp[30][21];
        stage0_col81[31] = pp[31][19];
        stage0_col82[0] = 1'b1;
        stage0_col82[1] = 1'b1;
        stage0_col82[2] = 1'b1;
        stage0_col82[3] = 1'b1;
        stage0_col82[4] = 1'b1;
        stage0_col82[5] = 1'b1;
        stage0_col82[6] = 1'b1;
        stage0_col82[7] = 1'b1;
        stage0_col82[8] = 1'b1;
        stage0_col82[9] = ~pp[9][64];
        stage0_col82[10] = 1'b1;
        stage0_col82[11] = pp[10][62];
        stage0_col82[12] = pp[11][60];
        stage0_col82[13] = pp[12][58];
        stage0_col82[14] = pp[13][56];
        stage0_col82[15] = pp[14][54];
        stage0_col82[16] = pp[15][52];
        stage0_col82[17] = pp[16][50];
        stage0_col82[18] = pp[17][48];
        stage0_col82[19] = pp[18][46];
        stage0_col82[20] = pp[19][44];
        stage0_col82[21] = pp[20][42];
        stage0_col82[22] = pp[21][40];
        stage0_col82[23] = pp[22][38];
        stage0_col82[24] = pp[23][36];
        stage0_col82[25] = pp[24][34];
        stage0_col82[26] = pp[25][32];
        stage0_col82[27] = pp[26][30];
        stage0_col82[28] = pp[27][28];
        stage0_col82[29] = pp[28][26];
        stage0_col82[30] = pp[29][24];
        stage0_col82[31] = pp[30][22];
        stage0_col82[32] = pp[31][20];
        stage0_col83[0] = 1'b1;
        stage0_col83[1] = 1'b1;
        stage0_col83[2] = 1'b1;
        stage0_col83[3] = 1'b1;
        stage0_col83[4] = 1'b1;
        stage0_col83[5] = 1'b1;
        stage0_col83[6] = 1'b1;
        stage0_col83[7] = 1'b1;
        stage0_col83[8] = 1'b1;
        stage0_col83[9] = 1'b1;
        stage0_col83[10] = pp[10][63];
        stage0_col83[11] = pp[11][61];
        stage0_col83[12] = pp[12][59];
        stage0_col83[13] = pp[13][57];
        stage0_col83[14] = pp[14][55];
        stage0_col83[15] = pp[15][53];
        stage0_col83[16] = pp[16][51];
        stage0_col83[17] = pp[17][49];
        stage0_col83[18] = pp[18][47];
        stage0_col83[19] = pp[19][45];
        stage0_col83[20] = pp[20][43];
        stage0_col83[21] = pp[21][41];
        stage0_col83[22] = pp[22][39];
        stage0_col83[23] = pp[23][37];
        stage0_col83[24] = pp[24][35];
        stage0_col83[25] = pp[25][33];
        stage0_col83[26] = pp[26][31];
        stage0_col83[27] = pp[27][29];
        stage0_col83[28] = pp[28][27];
        stage0_col83[29] = pp[29][25];
        stage0_col83[30] = pp[30][23];
        stage0_col83[31] = pp[31][21];
        stage0_col84[0] = 1'b1;
        stage0_col84[1] = 1'b1;
        stage0_col84[2] = 1'b1;
        stage0_col84[3] = 1'b1;
        stage0_col84[4] = 1'b1;
        stage0_col84[5] = 1'b1;
        stage0_col84[6] = 1'b1;
        stage0_col84[7] = 1'b1;
        stage0_col84[8] = 1'b1;
        stage0_col84[9] = 1'b1;
        stage0_col84[10] = ~pp[10][64];
        stage0_col84[11] = 1'b1;
        stage0_col84[12] = pp[11][62];
        stage0_col84[13] = pp[12][60];
        stage0_col84[14] = pp[13][58];
        stage0_col84[15] = pp[14][56];
        stage0_col84[16] = pp[15][54];
        stage0_col84[17] = pp[16][52];
        stage0_col84[18] = pp[17][50];
        stage0_col84[19] = pp[18][48];
        stage0_col84[20] = pp[19][46];
        stage0_col84[21] = pp[20][44];
        stage0_col84[22] = pp[21][42];
        stage0_col84[23] = pp[22][40];
        stage0_col84[24] = pp[23][38];
        stage0_col84[25] = pp[24][36];
        stage0_col84[26] = pp[25][34];
        stage0_col84[27] = pp[26][32];
        stage0_col84[28] = pp[27][30];
        stage0_col84[29] = pp[28][28];
        stage0_col84[30] = pp[29][26];
        stage0_col84[31] = pp[30][24];
        stage0_col84[32] = pp[31][22];
        stage0_col85[0] = 1'b1;
        stage0_col85[1] = 1'b1;
        stage0_col85[2] = 1'b1;
        stage0_col85[3] = 1'b1;
        stage0_col85[4] = 1'b1;
        stage0_col85[5] = 1'b1;
        stage0_col85[6] = 1'b1;
        stage0_col85[7] = 1'b1;
        stage0_col85[8] = 1'b1;
        stage0_col85[9] = 1'b1;
        stage0_col85[10] = 1'b1;
        stage0_col85[11] = pp[11][63];
        stage0_col85[12] = pp[12][61];
        stage0_col85[13] = pp[13][59];
        stage0_col85[14] = pp[14][57];
        stage0_col85[15] = pp[15][55];
        stage0_col85[16] = pp[16][53];
        stage0_col85[17] = pp[17][51];
        stage0_col85[18] = pp[18][49];
        stage0_col85[19] = pp[19][47];
        stage0_col85[20] = pp[20][45];
        stage0_col85[21] = pp[21][43];
        stage0_col85[22] = pp[22][41];
        stage0_col85[23] = pp[23][39];
        stage0_col85[24] = pp[24][37];
        stage0_col85[25] = pp[25][35];
        stage0_col85[26] = pp[26][33];
        stage0_col85[27] = pp[27][31];
        stage0_col85[28] = pp[28][29];
        stage0_col85[29] = pp[29][27];
        stage0_col85[30] = pp[30][25];
        stage0_col85[31] = pp[31][23];
        stage0_col86[0] = 1'b1;
        stage0_col86[1] = 1'b1;
        stage0_col86[2] = 1'b1;
        stage0_col86[3] = 1'b1;
        stage0_col86[4] = 1'b1;
        stage0_col86[5] = 1'b1;
        stage0_col86[6] = 1'b1;
        stage0_col86[7] = 1'b1;
        stage0_col86[8] = 1'b1;
        stage0_col86[9] = 1'b1;
        stage0_col86[10] = 1'b1;
        stage0_col86[11] = ~pp[11][64];
        stage0_col86[12] = 1'b1;
        stage0_col86[13] = pp[12][62];
        stage0_col86[14] = pp[13][60];
        stage0_col86[15] = pp[14][58];
        stage0_col86[16] = pp[15][56];
        stage0_col86[17] = pp[16][54];
        stage0_col86[18] = pp[17][52];
        stage0_col86[19] = pp[18][50];
        stage0_col86[20] = pp[19][48];
        stage0_col86[21] = pp[20][46];
        stage0_col86[22] = pp[21][44];
        stage0_col86[23] = pp[22][42];
        stage0_col86[24] = pp[23][40];
        stage0_col86[25] = pp[24][38];
        stage0_col86[26] = pp[25][36];
        stage0_col86[27] = pp[26][34];
        stage0_col86[28] = pp[27][32];
        stage0_col86[29] = pp[28][30];
        stage0_col86[30] = pp[29][28];
        stage0_col86[31] = pp[30][26];
        stage0_col86[32] = pp[31][24];
        stage0_col87[0] = 1'b1;
        stage0_col87[1] = 1'b1;
        stage0_col87[2] = 1'b1;
        stage0_col87[3] = 1'b1;
        stage0_col87[4] = 1'b1;
        stage0_col87[5] = 1'b1;
        stage0_col87[6] = 1'b1;
        stage0_col87[7] = 1'b1;
        stage0_col87[8] = 1'b1;
        stage0_col87[9] = 1'b1;
        stage0_col87[10] = 1'b1;
        stage0_col87[11] = 1'b1;
        stage0_col87[12] = pp[12][63];
        stage0_col87[13] = pp[13][61];
        stage0_col87[14] = pp[14][59];
        stage0_col87[15] = pp[15][57];
        stage0_col87[16] = pp[16][55];
        stage0_col87[17] = pp[17][53];
        stage0_col87[18] = pp[18][51];
        stage0_col87[19] = pp[19][49];
        stage0_col87[20] = pp[20][47];
        stage0_col87[21] = pp[21][45];
        stage0_col87[22] = pp[22][43];
        stage0_col87[23] = pp[23][41];
        stage0_col87[24] = pp[24][39];
        stage0_col87[25] = pp[25][37];
        stage0_col87[26] = pp[26][35];
        stage0_col87[27] = pp[27][33];
        stage0_col87[28] = pp[28][31];
        stage0_col87[29] = pp[29][29];
        stage0_col87[30] = pp[30][27];
        stage0_col87[31] = pp[31][25];
        stage0_col88[0] = 1'b1;
        stage0_col88[1] = 1'b1;
        stage0_col88[2] = 1'b1;
        stage0_col88[3] = 1'b1;
        stage0_col88[4] = 1'b1;
        stage0_col88[5] = 1'b1;
        stage0_col88[6] = 1'b1;
        stage0_col88[7] = 1'b1;
        stage0_col88[8] = 1'b1;
        stage0_col88[9] = 1'b1;
        stage0_col88[10] = 1'b1;
        stage0_col88[11] = 1'b1;
        stage0_col88[12] = ~pp[12][64];
        stage0_col88[13] = 1'b1;
        stage0_col88[14] = pp[13][62];
        stage0_col88[15] = pp[14][60];
        stage0_col88[16] = pp[15][58];
        stage0_col88[17] = pp[16][56];
        stage0_col88[18] = pp[17][54];
        stage0_col88[19] = pp[18][52];
        stage0_col88[20] = pp[19][50];
        stage0_col88[21] = pp[20][48];
        stage0_col88[22] = pp[21][46];
        stage0_col88[23] = pp[22][44];
        stage0_col88[24] = pp[23][42];
        stage0_col88[25] = pp[24][40];
        stage0_col88[26] = pp[25][38];
        stage0_col88[27] = pp[26][36];
        stage0_col88[28] = pp[27][34];
        stage0_col88[29] = pp[28][32];
        stage0_col88[30] = pp[29][30];
        stage0_col88[31] = pp[30][28];
        stage0_col88[32] = pp[31][26];
        stage0_col89[0] = 1'b1;
        stage0_col89[1] = 1'b1;
        stage0_col89[2] = 1'b1;
        stage0_col89[3] = 1'b1;
        stage0_col89[4] = 1'b1;
        stage0_col89[5] = 1'b1;
        stage0_col89[6] = 1'b1;
        stage0_col89[7] = 1'b1;
        stage0_col89[8] = 1'b1;
        stage0_col89[9] = 1'b1;
        stage0_col89[10] = 1'b1;
        stage0_col89[11] = 1'b1;
        stage0_col89[12] = 1'b1;
        stage0_col89[13] = pp[13][63];
        stage0_col89[14] = pp[14][61];
        stage0_col89[15] = pp[15][59];
        stage0_col89[16] = pp[16][57];
        stage0_col89[17] = pp[17][55];
        stage0_col89[18] = pp[18][53];
        stage0_col89[19] = pp[19][51];
        stage0_col89[20] = pp[20][49];
        stage0_col89[21] = pp[21][47];
        stage0_col89[22] = pp[22][45];
        stage0_col89[23] = pp[23][43];
        stage0_col89[24] = pp[24][41];
        stage0_col89[25] = pp[25][39];
        stage0_col89[26] = pp[26][37];
        stage0_col89[27] = pp[27][35];
        stage0_col89[28] = pp[28][33];
        stage0_col89[29] = pp[29][31];
        stage0_col89[30] = pp[30][29];
        stage0_col89[31] = pp[31][27];
        stage0_col90[0] = 1'b1;
        stage0_col90[1] = 1'b1;
        stage0_col90[2] = 1'b1;
        stage0_col90[3] = 1'b1;
        stage0_col90[4] = 1'b1;
        stage0_col90[5] = 1'b1;
        stage0_col90[6] = 1'b1;
        stage0_col90[7] = 1'b1;
        stage0_col90[8] = 1'b1;
        stage0_col90[9] = 1'b1;
        stage0_col90[10] = 1'b1;
        stage0_col90[11] = 1'b1;
        stage0_col90[12] = 1'b1;
        stage0_col90[13] = ~pp[13][64];
        stage0_col90[14] = 1'b1;
        stage0_col90[15] = pp[14][62];
        stage0_col90[16] = pp[15][60];
        stage0_col90[17] = pp[16][58];
        stage0_col90[18] = pp[17][56];
        stage0_col90[19] = pp[18][54];
        stage0_col90[20] = pp[19][52];
        stage0_col90[21] = pp[20][50];
        stage0_col90[22] = pp[21][48];
        stage0_col90[23] = pp[22][46];
        stage0_col90[24] = pp[23][44];
        stage0_col90[25] = pp[24][42];
        stage0_col90[26] = pp[25][40];
        stage0_col90[27] = pp[26][38];
        stage0_col90[28] = pp[27][36];
        stage0_col90[29] = pp[28][34];
        stage0_col90[30] = pp[29][32];
        stage0_col90[31] = pp[30][30];
        stage0_col90[32] = pp[31][28];
        stage0_col91[0] = 1'b1;
        stage0_col91[1] = 1'b1;
        stage0_col91[2] = 1'b1;
        stage0_col91[3] = 1'b1;
        stage0_col91[4] = 1'b1;
        stage0_col91[5] = 1'b1;
        stage0_col91[6] = 1'b1;
        stage0_col91[7] = 1'b1;
        stage0_col91[8] = 1'b1;
        stage0_col91[9] = 1'b1;
        stage0_col91[10] = 1'b1;
        stage0_col91[11] = 1'b1;
        stage0_col91[12] = 1'b1;
        stage0_col91[13] = 1'b1;
        stage0_col91[14] = pp[14][63];
        stage0_col91[15] = pp[15][61];
        stage0_col91[16] = pp[16][59];
        stage0_col91[17] = pp[17][57];
        stage0_col91[18] = pp[18][55];
        stage0_col91[19] = pp[19][53];
        stage0_col91[20] = pp[20][51];
        stage0_col91[21] = pp[21][49];
        stage0_col91[22] = pp[22][47];
        stage0_col91[23] = pp[23][45];
        stage0_col91[24] = pp[24][43];
        stage0_col91[25] = pp[25][41];
        stage0_col91[26] = pp[26][39];
        stage0_col91[27] = pp[27][37];
        stage0_col91[28] = pp[28][35];
        stage0_col91[29] = pp[29][33];
        stage0_col91[30] = pp[30][31];
        stage0_col91[31] = pp[31][29];
        stage0_col92[0] = 1'b1;
        stage0_col92[1] = 1'b1;
        stage0_col92[2] = 1'b1;
        stage0_col92[3] = 1'b1;
        stage0_col92[4] = 1'b1;
        stage0_col92[5] = 1'b1;
        stage0_col92[6] = 1'b1;
        stage0_col92[7] = 1'b1;
        stage0_col92[8] = 1'b1;
        stage0_col92[9] = 1'b1;
        stage0_col92[10] = 1'b1;
        stage0_col92[11] = 1'b1;
        stage0_col92[12] = 1'b1;
        stage0_col92[13] = 1'b1;
        stage0_col92[14] = ~pp[14][64];
        stage0_col92[15] = 1'b1;
        stage0_col92[16] = pp[15][62];
        stage0_col92[17] = pp[16][60];
        stage0_col92[18] = pp[17][58];
        stage0_col92[19] = pp[18][56];
        stage0_col92[20] = pp[19][54];
        stage0_col92[21] = pp[20][52];
        stage0_col92[22] = pp[21][50];
        stage0_col92[23] = pp[22][48];
        stage0_col92[24] = pp[23][46];
        stage0_col92[25] = pp[24][44];
        stage0_col92[26] = pp[25][42];
        stage0_col92[27] = pp[26][40];
        stage0_col92[28] = pp[27][38];
        stage0_col92[29] = pp[28][36];
        stage0_col92[30] = pp[29][34];
        stage0_col92[31] = pp[30][32];
        stage0_col92[32] = pp[31][30];
        stage0_col93[0] = 1'b1;
        stage0_col93[1] = 1'b1;
        stage0_col93[2] = 1'b1;
        stage0_col93[3] = 1'b1;
        stage0_col93[4] = 1'b1;
        stage0_col93[5] = 1'b1;
        stage0_col93[6] = 1'b1;
        stage0_col93[7] = 1'b1;
        stage0_col93[8] = 1'b1;
        stage0_col93[9] = 1'b1;
        stage0_col93[10] = 1'b1;
        stage0_col93[11] = 1'b1;
        stage0_col93[12] = 1'b1;
        stage0_col93[13] = 1'b1;
        stage0_col93[14] = 1'b1;
        stage0_col93[15] = pp[15][63];
        stage0_col93[16] = pp[16][61];
        stage0_col93[17] = pp[17][59];
        stage0_col93[18] = pp[18][57];
        stage0_col93[19] = pp[19][55];
        stage0_col93[20] = pp[20][53];
        stage0_col93[21] = pp[21][51];
        stage0_col93[22] = pp[22][49];
        stage0_col93[23] = pp[23][47];
        stage0_col93[24] = pp[24][45];
        stage0_col93[25] = pp[25][43];
        stage0_col93[26] = pp[26][41];
        stage0_col93[27] = pp[27][39];
        stage0_col93[28] = pp[28][37];
        stage0_col93[29] = pp[29][35];
        stage0_col93[30] = pp[30][33];
        stage0_col93[31] = pp[31][31];
        stage0_col94[0] = 1'b1;
        stage0_col94[1] = 1'b1;
        stage0_col94[2] = 1'b1;
        stage0_col94[3] = 1'b1;
        stage0_col94[4] = 1'b1;
        stage0_col94[5] = 1'b1;
        stage0_col94[6] = 1'b1;
        stage0_col94[7] = 1'b1;
        stage0_col94[8] = 1'b1;
        stage0_col94[9] = 1'b1;
        stage0_col94[10] = 1'b1;
        stage0_col94[11] = 1'b1;
        stage0_col94[12] = 1'b1;
        stage0_col94[13] = 1'b1;
        stage0_col94[14] = 1'b1;
        stage0_col94[15] = ~pp[15][64];
        stage0_col94[16] = 1'b1;
        stage0_col94[17] = pp[16][62];
        stage0_col94[18] = pp[17][60];
        stage0_col94[19] = pp[18][58];
        stage0_col94[20] = pp[19][56];
        stage0_col94[21] = pp[20][54];
        stage0_col94[22] = pp[21][52];
        stage0_col94[23] = pp[22][50];
        stage0_col94[24] = pp[23][48];
        stage0_col94[25] = pp[24][46];
        stage0_col94[26] = pp[25][44];
        stage0_col94[27] = pp[26][42];
        stage0_col94[28] = pp[27][40];
        stage0_col94[29] = pp[28][38];
        stage0_col94[30] = pp[29][36];
        stage0_col94[31] = pp[30][34];
        stage0_col94[32] = pp[31][32];
        stage0_col95[0] = 1'b1;
        stage0_col95[1] = 1'b1;
        stage0_col95[2] = 1'b1;
        stage0_col95[3] = 1'b1;
        stage0_col95[4] = 1'b1;
        stage0_col95[5] = 1'b1;
        stage0_col95[6] = 1'b1;
        stage0_col95[7] = 1'b1;
        stage0_col95[8] = 1'b1;
        stage0_col95[9] = 1'b1;
        stage0_col95[10] = 1'b1;
        stage0_col95[11] = 1'b1;
        stage0_col95[12] = 1'b1;
        stage0_col95[13] = 1'b1;
        stage0_col95[14] = 1'b1;
        stage0_col95[15] = 1'b1;
        stage0_col95[16] = pp[16][63];
        stage0_col95[17] = pp[17][61];
        stage0_col95[18] = pp[18][59];
        stage0_col95[19] = pp[19][57];
        stage0_col95[20] = pp[20][55];
        stage0_col95[21] = pp[21][53];
        stage0_col95[22] = pp[22][51];
        stage0_col95[23] = pp[23][49];
        stage0_col95[24] = pp[24][47];
        stage0_col95[25] = pp[25][45];
        stage0_col95[26] = pp[26][43];
        stage0_col95[27] = pp[27][41];
        stage0_col95[28] = pp[28][39];
        stage0_col95[29] = pp[29][37];
        stage0_col95[30] = pp[30][35];
        stage0_col95[31] = pp[31][33];
        stage0_col96[0] = 1'b1;
        stage0_col96[1] = 1'b1;
        stage0_col96[2] = 1'b1;
        stage0_col96[3] = 1'b1;
        stage0_col96[4] = 1'b1;
        stage0_col96[5] = 1'b1;
        stage0_col96[6] = 1'b1;
        stage0_col96[7] = 1'b1;
        stage0_col96[8] = 1'b1;
        stage0_col96[9] = 1'b1;
        stage0_col96[10] = 1'b1;
        stage0_col96[11] = 1'b1;
        stage0_col96[12] = 1'b1;
        stage0_col96[13] = 1'b1;
        stage0_col96[14] = 1'b1;
        stage0_col96[15] = 1'b1;
        stage0_col96[16] = ~pp[16][64];
        stage0_col96[17] = 1'b1;
        stage0_col96[18] = pp[17][62];
        stage0_col96[19] = pp[18][60];
        stage0_col96[20] = pp[19][58];
        stage0_col96[21] = pp[20][56];
        stage0_col96[22] = pp[21][54];
        stage0_col96[23] = pp[22][52];
        stage0_col96[24] = pp[23][50];
        stage0_col96[25] = pp[24][48];
        stage0_col96[26] = pp[25][46];
        stage0_col96[27] = pp[26][44];
        stage0_col96[28] = pp[27][42];
        stage0_col96[29] = pp[28][40];
        stage0_col96[30] = pp[29][38];
        stage0_col96[31] = pp[30][36];
        stage0_col96[32] = pp[31][34];
        stage0_col97[0] = 1'b1;
        stage0_col97[1] = 1'b1;
        stage0_col97[2] = 1'b1;
        stage0_col97[3] = 1'b1;
        stage0_col97[4] = 1'b1;
        stage0_col97[5] = 1'b1;
        stage0_col97[6] = 1'b1;
        stage0_col97[7] = 1'b1;
        stage0_col97[8] = 1'b1;
        stage0_col97[9] = 1'b1;
        stage0_col97[10] = 1'b1;
        stage0_col97[11] = 1'b1;
        stage0_col97[12] = 1'b1;
        stage0_col97[13] = 1'b1;
        stage0_col97[14] = 1'b1;
        stage0_col97[15] = 1'b1;
        stage0_col97[16] = 1'b1;
        stage0_col97[17] = pp[17][63];
        stage0_col97[18] = pp[18][61];
        stage0_col97[19] = pp[19][59];
        stage0_col97[20] = pp[20][57];
        stage0_col97[21] = pp[21][55];
        stage0_col97[22] = pp[22][53];
        stage0_col97[23] = pp[23][51];
        stage0_col97[24] = pp[24][49];
        stage0_col97[25] = pp[25][47];
        stage0_col97[26] = pp[26][45];
        stage0_col97[27] = pp[27][43];
        stage0_col97[28] = pp[28][41];
        stage0_col97[29] = pp[29][39];
        stage0_col97[30] = pp[30][37];
        stage0_col97[31] = pp[31][35];
        stage0_col98[0] = 1'b1;
        stage0_col98[1] = 1'b1;
        stage0_col98[2] = 1'b1;
        stage0_col98[3] = 1'b1;
        stage0_col98[4] = 1'b1;
        stage0_col98[5] = 1'b1;
        stage0_col98[6] = 1'b1;
        stage0_col98[7] = 1'b1;
        stage0_col98[8] = 1'b1;
        stage0_col98[9] = 1'b1;
        stage0_col98[10] = 1'b1;
        stage0_col98[11] = 1'b1;
        stage0_col98[12] = 1'b1;
        stage0_col98[13] = 1'b1;
        stage0_col98[14] = 1'b1;
        stage0_col98[15] = 1'b1;
        stage0_col98[16] = 1'b1;
        stage0_col98[17] = ~pp[17][64];
        stage0_col98[18] = 1'b1;
        stage0_col98[19] = pp[18][62];
        stage0_col98[20] = pp[19][60];
        stage0_col98[21] = pp[20][58];
        stage0_col98[22] = pp[21][56];
        stage0_col98[23] = pp[22][54];
        stage0_col98[24] = pp[23][52];
        stage0_col98[25] = pp[24][50];
        stage0_col98[26] = pp[25][48];
        stage0_col98[27] = pp[26][46];
        stage0_col98[28] = pp[27][44];
        stage0_col98[29] = pp[28][42];
        stage0_col98[30] = pp[29][40];
        stage0_col98[31] = pp[30][38];
        stage0_col98[32] = pp[31][36];
        stage0_col99[0] = 1'b1;
        stage0_col99[1] = 1'b1;
        stage0_col99[2] = 1'b1;
        stage0_col99[3] = 1'b1;
        stage0_col99[4] = 1'b1;
        stage0_col99[5] = 1'b1;
        stage0_col99[6] = 1'b1;
        stage0_col99[7] = 1'b1;
        stage0_col99[8] = 1'b1;
        stage0_col99[9] = 1'b1;
        stage0_col99[10] = 1'b1;
        stage0_col99[11] = 1'b1;
        stage0_col99[12] = 1'b1;
        stage0_col99[13] = 1'b1;
        stage0_col99[14] = 1'b1;
        stage0_col99[15] = 1'b1;
        stage0_col99[16] = 1'b1;
        stage0_col99[17] = 1'b1;
        stage0_col99[18] = pp[18][63];
        stage0_col99[19] = pp[19][61];
        stage0_col99[20] = pp[20][59];
        stage0_col99[21] = pp[21][57];
        stage0_col99[22] = pp[22][55];
        stage0_col99[23] = pp[23][53];
        stage0_col99[24] = pp[24][51];
        stage0_col99[25] = pp[25][49];
        stage0_col99[26] = pp[26][47];
        stage0_col99[27] = pp[27][45];
        stage0_col99[28] = pp[28][43];
        stage0_col99[29] = pp[29][41];
        stage0_col99[30] = pp[30][39];
        stage0_col99[31] = pp[31][37];
        stage0_col100[0] = 1'b1;
        stage0_col100[1] = 1'b1;
        stage0_col100[2] = 1'b1;
        stage0_col100[3] = 1'b1;
        stage0_col100[4] = 1'b1;
        stage0_col100[5] = 1'b1;
        stage0_col100[6] = 1'b1;
        stage0_col100[7] = 1'b1;
        stage0_col100[8] = 1'b1;
        stage0_col100[9] = 1'b1;
        stage0_col100[10] = 1'b1;
        stage0_col100[11] = 1'b1;
        stage0_col100[12] = 1'b1;
        stage0_col100[13] = 1'b1;
        stage0_col100[14] = 1'b1;
        stage0_col100[15] = 1'b1;
        stage0_col100[16] = 1'b1;
        stage0_col100[17] = 1'b1;
        stage0_col100[18] = ~pp[18][64];
        stage0_col100[19] = 1'b1;
        stage0_col100[20] = pp[19][62];
        stage0_col100[21] = pp[20][60];
        stage0_col100[22] = pp[21][58];
        stage0_col100[23] = pp[22][56];
        stage0_col100[24] = pp[23][54];
        stage0_col100[25] = pp[24][52];
        stage0_col100[26] = pp[25][50];
        stage0_col100[27] = pp[26][48];
        stage0_col100[28] = pp[27][46];
        stage0_col100[29] = pp[28][44];
        stage0_col100[30] = pp[29][42];
        stage0_col100[31] = pp[30][40];
        stage0_col100[32] = pp[31][38];
        stage0_col101[0] = 1'b1;
        stage0_col101[1] = 1'b1;
        stage0_col101[2] = 1'b1;
        stage0_col101[3] = 1'b1;
        stage0_col101[4] = 1'b1;
        stage0_col101[5] = 1'b1;
        stage0_col101[6] = 1'b1;
        stage0_col101[7] = 1'b1;
        stage0_col101[8] = 1'b1;
        stage0_col101[9] = 1'b1;
        stage0_col101[10] = 1'b1;
        stage0_col101[11] = 1'b1;
        stage0_col101[12] = 1'b1;
        stage0_col101[13] = 1'b1;
        stage0_col101[14] = 1'b1;
        stage0_col101[15] = 1'b1;
        stage0_col101[16] = 1'b1;
        stage0_col101[17] = 1'b1;
        stage0_col101[18] = 1'b1;
        stage0_col101[19] = pp[19][63];
        stage0_col101[20] = pp[20][61];
        stage0_col101[21] = pp[21][59];
        stage0_col101[22] = pp[22][57];
        stage0_col101[23] = pp[23][55];
        stage0_col101[24] = pp[24][53];
        stage0_col101[25] = pp[25][51];
        stage0_col101[26] = pp[26][49];
        stage0_col101[27] = pp[27][47];
        stage0_col101[28] = pp[28][45];
        stage0_col101[29] = pp[29][43];
        stage0_col101[30] = pp[30][41];
        stage0_col101[31] = pp[31][39];
        stage0_col102[0] = 1'b1;
        stage0_col102[1] = 1'b1;
        stage0_col102[2] = 1'b1;
        stage0_col102[3] = 1'b1;
        stage0_col102[4] = 1'b1;
        stage0_col102[5] = 1'b1;
        stage0_col102[6] = 1'b1;
        stage0_col102[7] = 1'b1;
        stage0_col102[8] = 1'b1;
        stage0_col102[9] = 1'b1;
        stage0_col102[10] = 1'b1;
        stage0_col102[11] = 1'b1;
        stage0_col102[12] = 1'b1;
        stage0_col102[13] = 1'b1;
        stage0_col102[14] = 1'b1;
        stage0_col102[15] = 1'b1;
        stage0_col102[16] = 1'b1;
        stage0_col102[17] = 1'b1;
        stage0_col102[18] = 1'b1;
        stage0_col102[19] = ~pp[19][64];
        stage0_col102[20] = 1'b1;
        stage0_col102[21] = pp[20][62];
        stage0_col102[22] = pp[21][60];
        stage0_col102[23] = pp[22][58];
        stage0_col102[24] = pp[23][56];
        stage0_col102[25] = pp[24][54];
        stage0_col102[26] = pp[25][52];
        stage0_col102[27] = pp[26][50];
        stage0_col102[28] = pp[27][48];
        stage0_col102[29] = pp[28][46];
        stage0_col102[30] = pp[29][44];
        stage0_col102[31] = pp[30][42];
        stage0_col102[32] = pp[31][40];
        stage0_col103[0] = 1'b1;
        stage0_col103[1] = 1'b1;
        stage0_col103[2] = 1'b1;
        stage0_col103[3] = 1'b1;
        stage0_col103[4] = 1'b1;
        stage0_col103[5] = 1'b1;
        stage0_col103[6] = 1'b1;
        stage0_col103[7] = 1'b1;
        stage0_col103[8] = 1'b1;
        stage0_col103[9] = 1'b1;
        stage0_col103[10] = 1'b1;
        stage0_col103[11] = 1'b1;
        stage0_col103[12] = 1'b1;
        stage0_col103[13] = 1'b1;
        stage0_col103[14] = 1'b1;
        stage0_col103[15] = 1'b1;
        stage0_col103[16] = 1'b1;
        stage0_col103[17] = 1'b1;
        stage0_col103[18] = 1'b1;
        stage0_col103[19] = 1'b1;
        stage0_col103[20] = pp[20][63];
        stage0_col103[21] = pp[21][61];
        stage0_col103[22] = pp[22][59];
        stage0_col103[23] = pp[23][57];
        stage0_col103[24] = pp[24][55];
        stage0_col103[25] = pp[25][53];
        stage0_col103[26] = pp[26][51];
        stage0_col103[27] = pp[27][49];
        stage0_col103[28] = pp[28][47];
        stage0_col103[29] = pp[29][45];
        stage0_col103[30] = pp[30][43];
        stage0_col103[31] = pp[31][41];
        stage0_col104[0] = 1'b1;
        stage0_col104[1] = 1'b1;
        stage0_col104[2] = 1'b1;
        stage0_col104[3] = 1'b1;
        stage0_col104[4] = 1'b1;
        stage0_col104[5] = 1'b1;
        stage0_col104[6] = 1'b1;
        stage0_col104[7] = 1'b1;
        stage0_col104[8] = 1'b1;
        stage0_col104[9] = 1'b1;
        stage0_col104[10] = 1'b1;
        stage0_col104[11] = 1'b1;
        stage0_col104[12] = 1'b1;
        stage0_col104[13] = 1'b1;
        stage0_col104[14] = 1'b1;
        stage0_col104[15] = 1'b1;
        stage0_col104[16] = 1'b1;
        stage0_col104[17] = 1'b1;
        stage0_col104[18] = 1'b1;
        stage0_col104[19] = 1'b1;
        stage0_col104[20] = ~pp[20][64];
        stage0_col104[21] = 1'b1;
        stage0_col104[22] = pp[21][62];
        stage0_col104[23] = pp[22][60];
        stage0_col104[24] = pp[23][58];
        stage0_col104[25] = pp[24][56];
        stage0_col104[26] = pp[25][54];
        stage0_col104[27] = pp[26][52];
        stage0_col104[28] = pp[27][50];
        stage0_col104[29] = pp[28][48];
        stage0_col104[30] = pp[29][46];
        stage0_col104[31] = pp[30][44];
        stage0_col104[32] = pp[31][42];
        stage0_col105[0] = 1'b1;
        stage0_col105[1] = 1'b1;
        stage0_col105[2] = 1'b1;
        stage0_col105[3] = 1'b1;
        stage0_col105[4] = 1'b1;
        stage0_col105[5] = 1'b1;
        stage0_col105[6] = 1'b1;
        stage0_col105[7] = 1'b1;
        stage0_col105[8] = 1'b1;
        stage0_col105[9] = 1'b1;
        stage0_col105[10] = 1'b1;
        stage0_col105[11] = 1'b1;
        stage0_col105[12] = 1'b1;
        stage0_col105[13] = 1'b1;
        stage0_col105[14] = 1'b1;
        stage0_col105[15] = 1'b1;
        stage0_col105[16] = 1'b1;
        stage0_col105[17] = 1'b1;
        stage0_col105[18] = 1'b1;
        stage0_col105[19] = 1'b1;
        stage0_col105[20] = 1'b1;
        stage0_col105[21] = pp[21][63];
        stage0_col105[22] = pp[22][61];
        stage0_col105[23] = pp[23][59];
        stage0_col105[24] = pp[24][57];
        stage0_col105[25] = pp[25][55];
        stage0_col105[26] = pp[26][53];
        stage0_col105[27] = pp[27][51];
        stage0_col105[28] = pp[28][49];
        stage0_col105[29] = pp[29][47];
        stage0_col105[30] = pp[30][45];
        stage0_col105[31] = pp[31][43];
        stage0_col106[0] = 1'b1;
        stage0_col106[1] = 1'b1;
        stage0_col106[2] = 1'b1;
        stage0_col106[3] = 1'b1;
        stage0_col106[4] = 1'b1;
        stage0_col106[5] = 1'b1;
        stage0_col106[6] = 1'b1;
        stage0_col106[7] = 1'b1;
        stage0_col106[8] = 1'b1;
        stage0_col106[9] = 1'b1;
        stage0_col106[10] = 1'b1;
        stage0_col106[11] = 1'b1;
        stage0_col106[12] = 1'b1;
        stage0_col106[13] = 1'b1;
        stage0_col106[14] = 1'b1;
        stage0_col106[15] = 1'b1;
        stage0_col106[16] = 1'b1;
        stage0_col106[17] = 1'b1;
        stage0_col106[18] = 1'b1;
        stage0_col106[19] = 1'b1;
        stage0_col106[20] = 1'b1;
        stage0_col106[21] = ~pp[21][64];
        stage0_col106[22] = 1'b1;
        stage0_col106[23] = pp[22][62];
        stage0_col106[24] = pp[23][60];
        stage0_col106[25] = pp[24][58];
        stage0_col106[26] = pp[25][56];
        stage0_col106[27] = pp[26][54];
        stage0_col106[28] = pp[27][52];
        stage0_col106[29] = pp[28][50];
        stage0_col106[30] = pp[29][48];
        stage0_col106[31] = pp[30][46];
        stage0_col106[32] = pp[31][44];
        stage0_col107[0] = 1'b1;
        stage0_col107[1] = 1'b1;
        stage0_col107[2] = 1'b1;
        stage0_col107[3] = 1'b1;
        stage0_col107[4] = 1'b1;
        stage0_col107[5] = 1'b1;
        stage0_col107[6] = 1'b1;
        stage0_col107[7] = 1'b1;
        stage0_col107[8] = 1'b1;
        stage0_col107[9] = 1'b1;
        stage0_col107[10] = 1'b1;
        stage0_col107[11] = 1'b1;
        stage0_col107[12] = 1'b1;
        stage0_col107[13] = 1'b1;
        stage0_col107[14] = 1'b1;
        stage0_col107[15] = 1'b1;
        stage0_col107[16] = 1'b1;
        stage0_col107[17] = 1'b1;
        stage0_col107[18] = 1'b1;
        stage0_col107[19] = 1'b1;
        stage0_col107[20] = 1'b1;
        stage0_col107[21] = 1'b1;
        stage0_col107[22] = pp[22][63];
        stage0_col107[23] = pp[23][61];
        stage0_col107[24] = pp[24][59];
        stage0_col107[25] = pp[25][57];
        stage0_col107[26] = pp[26][55];
        stage0_col107[27] = pp[27][53];
        stage0_col107[28] = pp[28][51];
        stage0_col107[29] = pp[29][49];
        stage0_col107[30] = pp[30][47];
        stage0_col107[31] = pp[31][45];
        stage0_col108[0] = 1'b1;
        stage0_col108[1] = 1'b1;
        stage0_col108[2] = 1'b1;
        stage0_col108[3] = 1'b1;
        stage0_col108[4] = 1'b1;
        stage0_col108[5] = 1'b1;
        stage0_col108[6] = 1'b1;
        stage0_col108[7] = 1'b1;
        stage0_col108[8] = 1'b1;
        stage0_col108[9] = 1'b1;
        stage0_col108[10] = 1'b1;
        stage0_col108[11] = 1'b1;
        stage0_col108[12] = 1'b1;
        stage0_col108[13] = 1'b1;
        stage0_col108[14] = 1'b1;
        stage0_col108[15] = 1'b1;
        stage0_col108[16] = 1'b1;
        stage0_col108[17] = 1'b1;
        stage0_col108[18] = 1'b1;
        stage0_col108[19] = 1'b1;
        stage0_col108[20] = 1'b1;
        stage0_col108[21] = 1'b1;
        stage0_col108[22] = ~pp[22][64];
        stage0_col108[23] = 1'b1;
        stage0_col108[24] = pp[23][62];
        stage0_col108[25] = pp[24][60];
        stage0_col108[26] = pp[25][58];
        stage0_col108[27] = pp[26][56];
        stage0_col108[28] = pp[27][54];
        stage0_col108[29] = pp[28][52];
        stage0_col108[30] = pp[29][50];
        stage0_col108[31] = pp[30][48];
        stage0_col108[32] = pp[31][46];
        stage0_col109[0] = 1'b1;
        stage0_col109[1] = 1'b1;
        stage0_col109[2] = 1'b1;
        stage0_col109[3] = 1'b1;
        stage0_col109[4] = 1'b1;
        stage0_col109[5] = 1'b1;
        stage0_col109[6] = 1'b1;
        stage0_col109[7] = 1'b1;
        stage0_col109[8] = 1'b1;
        stage0_col109[9] = 1'b1;
        stage0_col109[10] = 1'b1;
        stage0_col109[11] = 1'b1;
        stage0_col109[12] = 1'b1;
        stage0_col109[13] = 1'b1;
        stage0_col109[14] = 1'b1;
        stage0_col109[15] = 1'b1;
        stage0_col109[16] = 1'b1;
        stage0_col109[17] = 1'b1;
        stage0_col109[18] = 1'b1;
        stage0_col109[19] = 1'b1;
        stage0_col109[20] = 1'b1;
        stage0_col109[21] = 1'b1;
        stage0_col109[22] = 1'b1;
        stage0_col109[23] = pp[23][63];
        stage0_col109[24] = pp[24][61];
        stage0_col109[25] = pp[25][59];
        stage0_col109[26] = pp[26][57];
        stage0_col109[27] = pp[27][55];
        stage0_col109[28] = pp[28][53];
        stage0_col109[29] = pp[29][51];
        stage0_col109[30] = pp[30][49];
        stage0_col109[31] = pp[31][47];
        stage0_col110[0] = 1'b1;
        stage0_col110[1] = 1'b1;
        stage0_col110[2] = 1'b1;
        stage0_col110[3] = 1'b1;
        stage0_col110[4] = 1'b1;
        stage0_col110[5] = 1'b1;
        stage0_col110[6] = 1'b1;
        stage0_col110[7] = 1'b1;
        stage0_col110[8] = 1'b1;
        stage0_col110[9] = 1'b1;
        stage0_col110[10] = 1'b1;
        stage0_col110[11] = 1'b1;
        stage0_col110[12] = 1'b1;
        stage0_col110[13] = 1'b1;
        stage0_col110[14] = 1'b1;
        stage0_col110[15] = 1'b1;
        stage0_col110[16] = 1'b1;
        stage0_col110[17] = 1'b1;
        stage0_col110[18] = 1'b1;
        stage0_col110[19] = 1'b1;
        stage0_col110[20] = 1'b1;
        stage0_col110[21] = 1'b1;
        stage0_col110[22] = 1'b1;
        stage0_col110[23] = ~pp[23][64];
        stage0_col110[24] = 1'b1;
        stage0_col110[25] = pp[24][62];
        stage0_col110[26] = pp[25][60];
        stage0_col110[27] = pp[26][58];
        stage0_col110[28] = pp[27][56];
        stage0_col110[29] = pp[28][54];
        stage0_col110[30] = pp[29][52];
        stage0_col110[31] = pp[30][50];
        stage0_col110[32] = pp[31][48];
        stage0_col111[0] = 1'b1;
        stage0_col111[1] = 1'b1;
        stage0_col111[2] = 1'b1;
        stage0_col111[3] = 1'b1;
        stage0_col111[4] = 1'b1;
        stage0_col111[5] = 1'b1;
        stage0_col111[6] = 1'b1;
        stage0_col111[7] = 1'b1;
        stage0_col111[8] = 1'b1;
        stage0_col111[9] = 1'b1;
        stage0_col111[10] = 1'b1;
        stage0_col111[11] = 1'b1;
        stage0_col111[12] = 1'b1;
        stage0_col111[13] = 1'b1;
        stage0_col111[14] = 1'b1;
        stage0_col111[15] = 1'b1;
        stage0_col111[16] = 1'b1;
        stage0_col111[17] = 1'b1;
        stage0_col111[18] = 1'b1;
        stage0_col111[19] = 1'b1;
        stage0_col111[20] = 1'b1;
        stage0_col111[21] = 1'b1;
        stage0_col111[22] = 1'b1;
        stage0_col111[23] = 1'b1;
        stage0_col111[24] = pp[24][63];
        stage0_col111[25] = pp[25][61];
        stage0_col111[26] = pp[26][59];
        stage0_col111[27] = pp[27][57];
        stage0_col111[28] = pp[28][55];
        stage0_col111[29] = pp[29][53];
        stage0_col111[30] = pp[30][51];
        stage0_col111[31] = pp[31][49];
        stage0_col112[0] = 1'b1;
        stage0_col112[1] = 1'b1;
        stage0_col112[2] = 1'b1;
        stage0_col112[3] = 1'b1;
        stage0_col112[4] = 1'b1;
        stage0_col112[5] = 1'b1;
        stage0_col112[6] = 1'b1;
        stage0_col112[7] = 1'b1;
        stage0_col112[8] = 1'b1;
        stage0_col112[9] = 1'b1;
        stage0_col112[10] = 1'b1;
        stage0_col112[11] = 1'b1;
        stage0_col112[12] = 1'b1;
        stage0_col112[13] = 1'b1;
        stage0_col112[14] = 1'b1;
        stage0_col112[15] = 1'b1;
        stage0_col112[16] = 1'b1;
        stage0_col112[17] = 1'b1;
        stage0_col112[18] = 1'b1;
        stage0_col112[19] = 1'b1;
        stage0_col112[20] = 1'b1;
        stage0_col112[21] = 1'b1;
        stage0_col112[22] = 1'b1;
        stage0_col112[23] = 1'b1;
        stage0_col112[24] = ~pp[24][64];
        stage0_col112[25] = 1'b1;
        stage0_col112[26] = pp[25][62];
        stage0_col112[27] = pp[26][60];
        stage0_col112[28] = pp[27][58];
        stage0_col112[29] = pp[28][56];
        stage0_col112[30] = pp[29][54];
        stage0_col112[31] = pp[30][52];
        stage0_col112[32] = pp[31][50];
        stage0_col113[0] = 1'b1;
        stage0_col113[1] = 1'b1;
        stage0_col113[2] = 1'b1;
        stage0_col113[3] = 1'b1;
        stage0_col113[4] = 1'b1;
        stage0_col113[5] = 1'b1;
        stage0_col113[6] = 1'b1;
        stage0_col113[7] = 1'b1;
        stage0_col113[8] = 1'b1;
        stage0_col113[9] = 1'b1;
        stage0_col113[10] = 1'b1;
        stage0_col113[11] = 1'b1;
        stage0_col113[12] = 1'b1;
        stage0_col113[13] = 1'b1;
        stage0_col113[14] = 1'b1;
        stage0_col113[15] = 1'b1;
        stage0_col113[16] = 1'b1;
        stage0_col113[17] = 1'b1;
        stage0_col113[18] = 1'b1;
        stage0_col113[19] = 1'b1;
        stage0_col113[20] = 1'b1;
        stage0_col113[21] = 1'b1;
        stage0_col113[22] = 1'b1;
        stage0_col113[23] = 1'b1;
        stage0_col113[24] = 1'b1;
        stage0_col113[25] = pp[25][63];
        stage0_col113[26] = pp[26][61];
        stage0_col113[27] = pp[27][59];
        stage0_col113[28] = pp[28][57];
        stage0_col113[29] = pp[29][55];
        stage0_col113[30] = pp[30][53];
        stage0_col113[31] = pp[31][51];
        stage0_col114[0] = 1'b1;
        stage0_col114[1] = 1'b1;
        stage0_col114[2] = 1'b1;
        stage0_col114[3] = 1'b1;
        stage0_col114[4] = 1'b1;
        stage0_col114[5] = 1'b1;
        stage0_col114[6] = 1'b1;
        stage0_col114[7] = 1'b1;
        stage0_col114[8] = 1'b1;
        stage0_col114[9] = 1'b1;
        stage0_col114[10] = 1'b1;
        stage0_col114[11] = 1'b1;
        stage0_col114[12] = 1'b1;
        stage0_col114[13] = 1'b1;
        stage0_col114[14] = 1'b1;
        stage0_col114[15] = 1'b1;
        stage0_col114[16] = 1'b1;
        stage0_col114[17] = 1'b1;
        stage0_col114[18] = 1'b1;
        stage0_col114[19] = 1'b1;
        stage0_col114[20] = 1'b1;
        stage0_col114[21] = 1'b1;
        stage0_col114[22] = 1'b1;
        stage0_col114[23] = 1'b1;
        stage0_col114[24] = 1'b1;
        stage0_col114[25] = ~pp[25][64];
        stage0_col114[26] = 1'b1;
        stage0_col114[27] = pp[26][62];
        stage0_col114[28] = pp[27][60];
        stage0_col114[29] = pp[28][58];
        stage0_col114[30] = pp[29][56];
        stage0_col114[31] = pp[30][54];
        stage0_col114[32] = pp[31][52];
        stage0_col115[0] = 1'b1;
        stage0_col115[1] = 1'b1;
        stage0_col115[2] = 1'b1;
        stage0_col115[3] = 1'b1;
        stage0_col115[4] = 1'b1;
        stage0_col115[5] = 1'b1;
        stage0_col115[6] = 1'b1;
        stage0_col115[7] = 1'b1;
        stage0_col115[8] = 1'b1;
        stage0_col115[9] = 1'b1;
        stage0_col115[10] = 1'b1;
        stage0_col115[11] = 1'b1;
        stage0_col115[12] = 1'b1;
        stage0_col115[13] = 1'b1;
        stage0_col115[14] = 1'b1;
        stage0_col115[15] = 1'b1;
        stage0_col115[16] = 1'b1;
        stage0_col115[17] = 1'b1;
        stage0_col115[18] = 1'b1;
        stage0_col115[19] = 1'b1;
        stage0_col115[20] = 1'b1;
        stage0_col115[21] = 1'b1;
        stage0_col115[22] = 1'b1;
        stage0_col115[23] = 1'b1;
        stage0_col115[24] = 1'b1;
        stage0_col115[25] = 1'b1;
        stage0_col115[26] = pp[26][63];
        stage0_col115[27] = pp[27][61];
        stage0_col115[28] = pp[28][59];
        stage0_col115[29] = pp[29][57];
        stage0_col115[30] = pp[30][55];
        stage0_col115[31] = pp[31][53];
        stage0_col116[0] = 1'b1;
        stage0_col116[1] = 1'b1;
        stage0_col116[2] = 1'b1;
        stage0_col116[3] = 1'b1;
        stage0_col116[4] = 1'b1;
        stage0_col116[5] = 1'b1;
        stage0_col116[6] = 1'b1;
        stage0_col116[7] = 1'b1;
        stage0_col116[8] = 1'b1;
        stage0_col116[9] = 1'b1;
        stage0_col116[10] = 1'b1;
        stage0_col116[11] = 1'b1;
        stage0_col116[12] = 1'b1;
        stage0_col116[13] = 1'b1;
        stage0_col116[14] = 1'b1;
        stage0_col116[15] = 1'b1;
        stage0_col116[16] = 1'b1;
        stage0_col116[17] = 1'b1;
        stage0_col116[18] = 1'b1;
        stage0_col116[19] = 1'b1;
        stage0_col116[20] = 1'b1;
        stage0_col116[21] = 1'b1;
        stage0_col116[22] = 1'b1;
        stage0_col116[23] = 1'b1;
        stage0_col116[24] = 1'b1;
        stage0_col116[25] = 1'b1;
        stage0_col116[26] = ~pp[26][64];
        stage0_col116[27] = 1'b1;
        stage0_col116[28] = pp[27][62];
        stage0_col116[29] = pp[28][60];
        stage0_col116[30] = pp[29][58];
        stage0_col116[31] = pp[30][56];
        stage0_col116[32] = pp[31][54];
        stage0_col117[0] = 1'b1;
        stage0_col117[1] = 1'b1;
        stage0_col117[2] = 1'b1;
        stage0_col117[3] = 1'b1;
        stage0_col117[4] = 1'b1;
        stage0_col117[5] = 1'b1;
        stage0_col117[6] = 1'b1;
        stage0_col117[7] = 1'b1;
        stage0_col117[8] = 1'b1;
        stage0_col117[9] = 1'b1;
        stage0_col117[10] = 1'b1;
        stage0_col117[11] = 1'b1;
        stage0_col117[12] = 1'b1;
        stage0_col117[13] = 1'b1;
        stage0_col117[14] = 1'b1;
        stage0_col117[15] = 1'b1;
        stage0_col117[16] = 1'b1;
        stage0_col117[17] = 1'b1;
        stage0_col117[18] = 1'b1;
        stage0_col117[19] = 1'b1;
        stage0_col117[20] = 1'b1;
        stage0_col117[21] = 1'b1;
        stage0_col117[22] = 1'b1;
        stage0_col117[23] = 1'b1;
        stage0_col117[24] = 1'b1;
        stage0_col117[25] = 1'b1;
        stage0_col117[26] = 1'b1;
        stage0_col117[27] = pp[27][63];
        stage0_col117[28] = pp[28][61];
        stage0_col117[29] = pp[29][59];
        stage0_col117[30] = pp[30][57];
        stage0_col117[31] = pp[31][55];
        stage0_col118[0] = 1'b1;
        stage0_col118[1] = 1'b1;
        stage0_col118[2] = 1'b1;
        stage0_col118[3] = 1'b1;
        stage0_col118[4] = 1'b1;
        stage0_col118[5] = 1'b1;
        stage0_col118[6] = 1'b1;
        stage0_col118[7] = 1'b1;
        stage0_col118[8] = 1'b1;
        stage0_col118[9] = 1'b1;
        stage0_col118[10] = 1'b1;
        stage0_col118[11] = 1'b1;
        stage0_col118[12] = 1'b1;
        stage0_col118[13] = 1'b1;
        stage0_col118[14] = 1'b1;
        stage0_col118[15] = 1'b1;
        stage0_col118[16] = 1'b1;
        stage0_col118[17] = 1'b1;
        stage0_col118[18] = 1'b1;
        stage0_col118[19] = 1'b1;
        stage0_col118[20] = 1'b1;
        stage0_col118[21] = 1'b1;
        stage0_col118[22] = 1'b1;
        stage0_col118[23] = 1'b1;
        stage0_col118[24] = 1'b1;
        stage0_col118[25] = 1'b1;
        stage0_col118[26] = 1'b1;
        stage0_col118[27] = ~pp[27][64];
        stage0_col118[28] = 1'b1;
        stage0_col118[29] = pp[28][62];
        stage0_col118[30] = pp[29][60];
        stage0_col118[31] = pp[30][58];
        stage0_col118[32] = pp[31][56];
        stage0_col119[0] = 1'b1;
        stage0_col119[1] = 1'b1;
        stage0_col119[2] = 1'b1;
        stage0_col119[3] = 1'b1;
        stage0_col119[4] = 1'b1;
        stage0_col119[5] = 1'b1;
        stage0_col119[6] = 1'b1;
        stage0_col119[7] = 1'b1;
        stage0_col119[8] = 1'b1;
        stage0_col119[9] = 1'b1;
        stage0_col119[10] = 1'b1;
        stage0_col119[11] = 1'b1;
        stage0_col119[12] = 1'b1;
        stage0_col119[13] = 1'b1;
        stage0_col119[14] = 1'b1;
        stage0_col119[15] = 1'b1;
        stage0_col119[16] = 1'b1;
        stage0_col119[17] = 1'b1;
        stage0_col119[18] = 1'b1;
        stage0_col119[19] = 1'b1;
        stage0_col119[20] = 1'b1;
        stage0_col119[21] = 1'b1;
        stage0_col119[22] = 1'b1;
        stage0_col119[23] = 1'b1;
        stage0_col119[24] = 1'b1;
        stage0_col119[25] = 1'b1;
        stage0_col119[26] = 1'b1;
        stage0_col119[27] = 1'b1;
        stage0_col119[28] = pp[28][63];
        stage0_col119[29] = pp[29][61];
        stage0_col119[30] = pp[30][59];
        stage0_col119[31] = pp[31][57];
        stage0_col120[0] = 1'b1;
        stage0_col120[1] = 1'b1;
        stage0_col120[2] = 1'b1;
        stage0_col120[3] = 1'b1;
        stage0_col120[4] = 1'b1;
        stage0_col120[5] = 1'b1;
        stage0_col120[6] = 1'b1;
        stage0_col120[7] = 1'b1;
        stage0_col120[8] = 1'b1;
        stage0_col120[9] = 1'b1;
        stage0_col120[10] = 1'b1;
        stage0_col120[11] = 1'b1;
        stage0_col120[12] = 1'b1;
        stage0_col120[13] = 1'b1;
        stage0_col120[14] = 1'b1;
        stage0_col120[15] = 1'b1;
        stage0_col120[16] = 1'b1;
        stage0_col120[17] = 1'b1;
        stage0_col120[18] = 1'b1;
        stage0_col120[19] = 1'b1;
        stage0_col120[20] = 1'b1;
        stage0_col120[21] = 1'b1;
        stage0_col120[22] = 1'b1;
        stage0_col120[23] = 1'b1;
        stage0_col120[24] = 1'b1;
        stage0_col120[25] = 1'b1;
        stage0_col120[26] = 1'b1;
        stage0_col120[27] = 1'b1;
        stage0_col120[28] = ~pp[28][64];
        stage0_col120[29] = 1'b1;
        stage0_col120[30] = pp[29][62];
        stage0_col120[31] = pp[30][60];
        stage0_col120[32] = pp[31][58];
        stage0_col121[0] = 1'b1;
        stage0_col121[1] = 1'b1;
        stage0_col121[2] = 1'b1;
        stage0_col121[3] = 1'b1;
        stage0_col121[4] = 1'b1;
        stage0_col121[5] = 1'b1;
        stage0_col121[6] = 1'b1;
        stage0_col121[7] = 1'b1;
        stage0_col121[8] = 1'b1;
        stage0_col121[9] = 1'b1;
        stage0_col121[10] = 1'b1;
        stage0_col121[11] = 1'b1;
        stage0_col121[12] = 1'b1;
        stage0_col121[13] = 1'b1;
        stage0_col121[14] = 1'b1;
        stage0_col121[15] = 1'b1;
        stage0_col121[16] = 1'b1;
        stage0_col121[17] = 1'b1;
        stage0_col121[18] = 1'b1;
        stage0_col121[19] = 1'b1;
        stage0_col121[20] = 1'b1;
        stage0_col121[21] = 1'b1;
        stage0_col121[22] = 1'b1;
        stage0_col121[23] = 1'b1;
        stage0_col121[24] = 1'b1;
        stage0_col121[25] = 1'b1;
        stage0_col121[26] = 1'b1;
        stage0_col121[27] = 1'b1;
        stage0_col121[28] = 1'b1;
        stage0_col121[29] = pp[29][63];
        stage0_col121[30] = pp[30][61];
        stage0_col121[31] = pp[31][59];
        stage0_col122[0] = 1'b1;
        stage0_col122[1] = 1'b1;
        stage0_col122[2] = 1'b1;
        stage0_col122[3] = 1'b1;
        stage0_col122[4] = 1'b1;
        stage0_col122[5] = 1'b1;
        stage0_col122[6] = 1'b1;
        stage0_col122[7] = 1'b1;
        stage0_col122[8] = 1'b1;
        stage0_col122[9] = 1'b1;
        stage0_col122[10] = 1'b1;
        stage0_col122[11] = 1'b1;
        stage0_col122[12] = 1'b1;
        stage0_col122[13] = 1'b1;
        stage0_col122[14] = 1'b1;
        stage0_col122[15] = 1'b1;
        stage0_col122[16] = 1'b1;
        stage0_col122[17] = 1'b1;
        stage0_col122[18] = 1'b1;
        stage0_col122[19] = 1'b1;
        stage0_col122[20] = 1'b1;
        stage0_col122[21] = 1'b1;
        stage0_col122[22] = 1'b1;
        stage0_col122[23] = 1'b1;
        stage0_col122[24] = 1'b1;
        stage0_col122[25] = 1'b1;
        stage0_col122[26] = 1'b1;
        stage0_col122[27] = 1'b1;
        stage0_col122[28] = 1'b1;
        stage0_col122[29] = ~pp[29][64];
        stage0_col122[30] = 1'b1;
        stage0_col122[31] = pp[30][62];
        stage0_col122[32] = pp[31][60];
        stage0_col123[0] = 1'b1;
        stage0_col123[1] = 1'b1;
        stage0_col123[2] = 1'b1;
        stage0_col123[3] = 1'b1;
        stage0_col123[4] = 1'b1;
        stage0_col123[5] = 1'b1;
        stage0_col123[6] = 1'b1;
        stage0_col123[7] = 1'b1;
        stage0_col123[8] = 1'b1;
        stage0_col123[9] = 1'b1;
        stage0_col123[10] = 1'b1;
        stage0_col123[11] = 1'b1;
        stage0_col123[12] = 1'b1;
        stage0_col123[13] = 1'b1;
        stage0_col123[14] = 1'b1;
        stage0_col123[15] = 1'b1;
        stage0_col123[16] = 1'b1;
        stage0_col123[17] = 1'b1;
        stage0_col123[18] = 1'b1;
        stage0_col123[19] = 1'b1;
        stage0_col123[20] = 1'b1;
        stage0_col123[21] = 1'b1;
        stage0_col123[22] = 1'b1;
        stage0_col123[23] = 1'b1;
        stage0_col123[24] = 1'b1;
        stage0_col123[25] = 1'b1;
        stage0_col123[26] = 1'b1;
        stage0_col123[27] = 1'b1;
        stage0_col123[28] = 1'b1;
        stage0_col123[29] = 1'b1;
        stage0_col123[30] = pp[30][63];
        stage0_col123[31] = pp[31][61];
        stage0_col124[0] = 1'b1;
        stage0_col124[1] = 1'b1;
        stage0_col124[2] = 1'b1;
        stage0_col124[3] = 1'b1;
        stage0_col124[4] = 1'b1;
        stage0_col124[5] = 1'b1;
        stage0_col124[6] = 1'b1;
        stage0_col124[7] = 1'b1;
        stage0_col124[8] = 1'b1;
        stage0_col124[9] = 1'b1;
        stage0_col124[10] = 1'b1;
        stage0_col124[11] = 1'b1;
        stage0_col124[12] = 1'b1;
        stage0_col124[13] = 1'b1;
        stage0_col124[14] = 1'b1;
        stage0_col124[15] = 1'b1;
        stage0_col124[16] = 1'b1;
        stage0_col124[17] = 1'b1;
        stage0_col124[18] = 1'b1;
        stage0_col124[19] = 1'b1;
        stage0_col124[20] = 1'b1;
        stage0_col124[21] = 1'b1;
        stage0_col124[22] = 1'b1;
        stage0_col124[23] = 1'b1;
        stage0_col124[24] = 1'b1;
        stage0_col124[25] = 1'b1;
        stage0_col124[26] = 1'b1;
        stage0_col124[27] = 1'b1;
        stage0_col124[28] = 1'b1;
        stage0_col124[29] = 1'b1;
        stage0_col124[30] = ~pp[30][64];
        stage0_col124[31] = 1'b1;
        stage0_col124[32] = pp[31][62];
        stage0_col125[0] = 1'b1;
        stage0_col125[1] = 1'b1;
        stage0_col125[2] = 1'b1;
        stage0_col125[3] = 1'b1;
        stage0_col125[4] = 1'b1;
        stage0_col125[5] = 1'b1;
        stage0_col125[6] = 1'b1;
        stage0_col125[7] = 1'b1;
        stage0_col125[8] = 1'b1;
        stage0_col125[9] = 1'b1;
        stage0_col125[10] = 1'b1;
        stage0_col125[11] = 1'b1;
        stage0_col125[12] = 1'b1;
        stage0_col125[13] = 1'b1;
        stage0_col125[14] = 1'b1;
        stage0_col125[15] = 1'b1;
        stage0_col125[16] = 1'b1;
        stage0_col125[17] = 1'b1;
        stage0_col125[18] = 1'b1;
        stage0_col125[19] = 1'b1;
        stage0_col125[20] = 1'b1;
        stage0_col125[21] = 1'b1;
        stage0_col125[22] = 1'b1;
        stage0_col125[23] = 1'b1;
        stage0_col125[24] = 1'b1;
        stage0_col125[25] = 1'b1;
        stage0_col125[26] = 1'b1;
        stage0_col125[27] = 1'b1;
        stage0_col125[28] = 1'b1;
        stage0_col125[29] = 1'b1;
        stage0_col125[30] = 1'b1;
        stage0_col125[31] = pp[31][63];
        stage0_col126[0] = 1'b1;
        stage0_col126[1] = 1'b1;
        stage0_col126[2] = 1'b1;
        stage0_col126[3] = 1'b1;
        stage0_col126[4] = 1'b1;
        stage0_col126[5] = 1'b1;
        stage0_col126[6] = 1'b1;
        stage0_col126[7] = 1'b1;
        stage0_col126[8] = 1'b1;
        stage0_col126[9] = 1'b1;
        stage0_col126[10] = 1'b1;
        stage0_col126[11] = 1'b1;
        stage0_col126[12] = 1'b1;
        stage0_col126[13] = 1'b1;
        stage0_col126[14] = 1'b1;
        stage0_col126[15] = 1'b1;
        stage0_col126[16] = 1'b1;
        stage0_col126[17] = 1'b1;
        stage0_col126[18] = 1'b1;
        stage0_col126[19] = 1'b1;
        stage0_col126[20] = 1'b1;
        stage0_col126[21] = 1'b1;
        stage0_col126[22] = 1'b1;
        stage0_col126[23] = 1'b1;
        stage0_col126[24] = 1'b1;
        stage0_col126[25] = 1'b1;
        stage0_col126[26] = 1'b1;
        stage0_col126[27] = 1'b1;
        stage0_col126[28] = 1'b1;
        stage0_col126[29] = 1'b1;
        stage0_col126[30] = 1'b1;
        stage0_col126[31] = ~pp[31][64];
        stage0_col126[32] = 1'b1;
        stage0_col127[0] = 1'b1;
        stage0_col127[1] = 1'b1;
        stage0_col127[2] = 1'b1;
        stage0_col127[3] = 1'b1;
        stage0_col127[4] = 1'b1;
        stage0_col127[5] = 1'b1;
        stage0_col127[6] = 1'b1;
        stage0_col127[7] = 1'b1;
        stage0_col127[8] = 1'b1;
        stage0_col127[9] = 1'b1;
        stage0_col127[10] = 1'b1;
        stage0_col127[11] = 1'b1;
        stage0_col127[12] = 1'b1;
        stage0_col127[13] = 1'b1;
        stage0_col127[14] = 1'b1;
        stage0_col127[15] = 1'b1;
        stage0_col127[16] = 1'b1;
        stage0_col127[17] = 1'b1;
        stage0_col127[18] = 1'b1;
        stage0_col127[19] = 1'b1;
        stage0_col127[20] = 1'b1;
        stage0_col127[21] = 1'b1;
        stage0_col127[22] = 1'b1;
        stage0_col127[23] = 1'b1;
        stage0_col127[24] = 1'b1;
        stage0_col127[25] = 1'b1;
        stage0_col127[26] = 1'b1;
        stage0_col127[27] = 1'b1;
        stage0_col127[28] = 1'b1;
        stage0_col127[29] = 1'b1;
        stage0_col127[30] = 1'b1;
        stage0_col127[31] = 1'b1;
    end


    // Stage 1: Reduction
    fa fa_s0_c2_n0 (
        .a(stage0_col2[0]),
        .b(stage0_col2[1]),
        .c_in(stage0_col2[2]),
        .s(fa_s0_c2_n0_s),
        .c_out(fa_s0_c2_n0_c)
    );

    fa fa_s0_c4_n1 (
        .a(stage0_col4[0]),
        .b(stage0_col4[1]),
        .c_in(stage0_col4[2]),
        .s(fa_s0_c4_n1_s),
        .c_out(fa_s0_c4_n1_c)
    );

    fa fa_s0_c5_n2 (
        .a(stage0_col5[0]),
        .b(stage0_col5[1]),
        .c_in(stage0_col5[2]),
        .s(fa_s0_c5_n2_s),
        .c_out(fa_s0_c5_n2_c)
    );

    fa fa_s0_c6_n3 (
        .a(stage0_col6[0]),
        .b(stage0_col6[1]),
        .c_in(stage0_col6[2]),
        .s(fa_s0_c6_n3_s),
        .c_out(fa_s0_c6_n3_c)
    );

    fa fa_s0_c7_n4 (
        .a(stage0_col7[0]),
        .b(stage0_col7[1]),
        .c_in(stage0_col7[2]),
        .s(fa_s0_c7_n4_s),
        .c_out(fa_s0_c7_n4_c)
    );

    fa fa_s0_c8_n5 (
        .a(stage0_col8[0]),
        .b(stage0_col8[1]),
        .c_in(stage0_col8[2]),
        .s(fa_s0_c8_n5_s),
        .c_out(fa_s0_c8_n5_c)
    );

    fa fa_s0_c8_n6 (
        .a(stage0_col8[3]),
        .b(stage0_col8[4]),
        .c_in(stage0_col8[5]),
        .s(fa_s0_c8_n6_s),
        .c_out(fa_s0_c8_n6_c)
    );

    fa fa_s0_c9_n7 (
        .a(stage0_col9[0]),
        .b(stage0_col9[1]),
        .c_in(stage0_col9[2]),
        .s(fa_s0_c9_n7_s),
        .c_out(fa_s0_c9_n7_c)
    );

    fa fa_s0_c10_n8 (
        .a(stage0_col10[0]),
        .b(stage0_col10[1]),
        .c_in(stage0_col10[2]),
        .s(fa_s0_c10_n8_s),
        .c_out(fa_s0_c10_n8_c)
    );

    fa fa_s0_c10_n9 (
        .a(stage0_col10[3]),
        .b(stage0_col10[4]),
        .c_in(stage0_col10[5]),
        .s(fa_s0_c10_n9_s),
        .c_out(fa_s0_c10_n9_c)
    );

    fa fa_s0_c11_n10 (
        .a(stage0_col11[0]),
        .b(stage0_col11[1]),
        .c_in(stage0_col11[2]),
        .s(fa_s0_c11_n10_s),
        .c_out(fa_s0_c11_n10_c)
    );

    fa fa_s0_c11_n11 (
        .a(stage0_col11[3]),
        .b(stage0_col11[4]),
        .c_in(stage0_col11[5]),
        .s(fa_s0_c11_n11_s),
        .c_out(fa_s0_c11_n11_c)
    );

    fa fa_s0_c12_n12 (
        .a(stage0_col12[0]),
        .b(stage0_col12[1]),
        .c_in(stage0_col12[2]),
        .s(fa_s0_c12_n12_s),
        .c_out(fa_s0_c12_n12_c)
    );

    fa fa_s0_c12_n13 (
        .a(stage0_col12[3]),
        .b(stage0_col12[4]),
        .c_in(stage0_col12[5]),
        .s(fa_s0_c12_n13_s),
        .c_out(fa_s0_c12_n13_c)
    );

    fa fa_s0_c13_n14 (
        .a(stage0_col13[0]),
        .b(stage0_col13[1]),
        .c_in(stage0_col13[2]),
        .s(fa_s0_c13_n14_s),
        .c_out(fa_s0_c13_n14_c)
    );

    fa fa_s0_c13_n15 (
        .a(stage0_col13[3]),
        .b(stage0_col13[4]),
        .c_in(stage0_col13[5]),
        .s(fa_s0_c13_n15_s),
        .c_out(fa_s0_c13_n15_c)
    );

    fa fa_s0_c14_n16 (
        .a(stage0_col14[0]),
        .b(stage0_col14[1]),
        .c_in(stage0_col14[2]),
        .s(fa_s0_c14_n16_s),
        .c_out(fa_s0_c14_n16_c)
    );

    fa fa_s0_c14_n17 (
        .a(stage0_col14[3]),
        .b(stage0_col14[4]),
        .c_in(stage0_col14[5]),
        .s(fa_s0_c14_n17_s),
        .c_out(fa_s0_c14_n17_c)
    );

    fa fa_s0_c14_n18 (
        .a(stage0_col14[6]),
        .b(stage0_col14[7]),
        .c_in(stage0_col14[8]),
        .s(fa_s0_c14_n18_s),
        .c_out(fa_s0_c14_n18_c)
    );

    fa fa_s0_c15_n19 (
        .a(stage0_col15[0]),
        .b(stage0_col15[1]),
        .c_in(stage0_col15[2]),
        .s(fa_s0_c15_n19_s),
        .c_out(fa_s0_c15_n19_c)
    );

    fa fa_s0_c15_n20 (
        .a(stage0_col15[3]),
        .b(stage0_col15[4]),
        .c_in(stage0_col15[5]),
        .s(fa_s0_c15_n20_s),
        .c_out(fa_s0_c15_n20_c)
    );

    fa fa_s0_c16_n21 (
        .a(stage0_col16[0]),
        .b(stage0_col16[1]),
        .c_in(stage0_col16[2]),
        .s(fa_s0_c16_n21_s),
        .c_out(fa_s0_c16_n21_c)
    );

    fa fa_s0_c16_n22 (
        .a(stage0_col16[3]),
        .b(stage0_col16[4]),
        .c_in(stage0_col16[5]),
        .s(fa_s0_c16_n22_s),
        .c_out(fa_s0_c16_n22_c)
    );

    fa fa_s0_c16_n23 (
        .a(stage0_col16[6]),
        .b(stage0_col16[7]),
        .c_in(stage0_col16[8]),
        .s(fa_s0_c16_n23_s),
        .c_out(fa_s0_c16_n23_c)
    );

    fa fa_s0_c17_n24 (
        .a(stage0_col17[0]),
        .b(stage0_col17[1]),
        .c_in(stage0_col17[2]),
        .s(fa_s0_c17_n24_s),
        .c_out(fa_s0_c17_n24_c)
    );

    fa fa_s0_c17_n25 (
        .a(stage0_col17[3]),
        .b(stage0_col17[4]),
        .c_in(stage0_col17[5]),
        .s(fa_s0_c17_n25_s),
        .c_out(fa_s0_c17_n25_c)
    );

    fa fa_s0_c17_n26 (
        .a(stage0_col17[6]),
        .b(stage0_col17[7]),
        .c_in(stage0_col17[8]),
        .s(fa_s0_c17_n26_s),
        .c_out(fa_s0_c17_n26_c)
    );

    fa fa_s0_c18_n27 (
        .a(stage0_col18[0]),
        .b(stage0_col18[1]),
        .c_in(stage0_col18[2]),
        .s(fa_s0_c18_n27_s),
        .c_out(fa_s0_c18_n27_c)
    );

    fa fa_s0_c18_n28 (
        .a(stage0_col18[3]),
        .b(stage0_col18[4]),
        .c_in(stage0_col18[5]),
        .s(fa_s0_c18_n28_s),
        .c_out(fa_s0_c18_n28_c)
    );

    fa fa_s0_c18_n29 (
        .a(stage0_col18[6]),
        .b(stage0_col18[7]),
        .c_in(stage0_col18[8]),
        .s(fa_s0_c18_n29_s),
        .c_out(fa_s0_c18_n29_c)
    );

    fa fa_s0_c19_n30 (
        .a(stage0_col19[0]),
        .b(stage0_col19[1]),
        .c_in(stage0_col19[2]),
        .s(fa_s0_c19_n30_s),
        .c_out(fa_s0_c19_n30_c)
    );

    fa fa_s0_c19_n31 (
        .a(stage0_col19[3]),
        .b(stage0_col19[4]),
        .c_in(stage0_col19[5]),
        .s(fa_s0_c19_n31_s),
        .c_out(fa_s0_c19_n31_c)
    );

    fa fa_s0_c19_n32 (
        .a(stage0_col19[6]),
        .b(stage0_col19[7]),
        .c_in(stage0_col19[8]),
        .s(fa_s0_c19_n32_s),
        .c_out(fa_s0_c19_n32_c)
    );

    fa fa_s0_c20_n33 (
        .a(stage0_col20[0]),
        .b(stage0_col20[1]),
        .c_in(stage0_col20[2]),
        .s(fa_s0_c20_n33_s),
        .c_out(fa_s0_c20_n33_c)
    );

    fa fa_s0_c20_n34 (
        .a(stage0_col20[3]),
        .b(stage0_col20[4]),
        .c_in(stage0_col20[5]),
        .s(fa_s0_c20_n34_s),
        .c_out(fa_s0_c20_n34_c)
    );

    fa fa_s0_c20_n35 (
        .a(stage0_col20[6]),
        .b(stage0_col20[7]),
        .c_in(stage0_col20[8]),
        .s(fa_s0_c20_n35_s),
        .c_out(fa_s0_c20_n35_c)
    );

    fa fa_s0_c20_n36 (
        .a(stage0_col20[9]),
        .b(stage0_col20[10]),
        .c_in(stage0_col20[11]),
        .s(fa_s0_c20_n36_s),
        .c_out(fa_s0_c20_n36_c)
    );

    fa fa_s0_c21_n37 (
        .a(stage0_col21[0]),
        .b(stage0_col21[1]),
        .c_in(stage0_col21[2]),
        .s(fa_s0_c21_n37_s),
        .c_out(fa_s0_c21_n37_c)
    );

    fa fa_s0_c21_n38 (
        .a(stage0_col21[3]),
        .b(stage0_col21[4]),
        .c_in(stage0_col21[5]),
        .s(fa_s0_c21_n38_s),
        .c_out(fa_s0_c21_n38_c)
    );

    fa fa_s0_c21_n39 (
        .a(stage0_col21[6]),
        .b(stage0_col21[7]),
        .c_in(stage0_col21[8]),
        .s(fa_s0_c21_n39_s),
        .c_out(fa_s0_c21_n39_c)
    );

    fa fa_s0_c22_n40 (
        .a(stage0_col22[0]),
        .b(stage0_col22[1]),
        .c_in(stage0_col22[2]),
        .s(fa_s0_c22_n40_s),
        .c_out(fa_s0_c22_n40_c)
    );

    fa fa_s0_c22_n41 (
        .a(stage0_col22[3]),
        .b(stage0_col22[4]),
        .c_in(stage0_col22[5]),
        .s(fa_s0_c22_n41_s),
        .c_out(fa_s0_c22_n41_c)
    );

    fa fa_s0_c22_n42 (
        .a(stage0_col22[6]),
        .b(stage0_col22[7]),
        .c_in(stage0_col22[8]),
        .s(fa_s0_c22_n42_s),
        .c_out(fa_s0_c22_n42_c)
    );

    fa fa_s0_c22_n43 (
        .a(stage0_col22[9]),
        .b(stage0_col22[10]),
        .c_in(stage0_col22[11]),
        .s(fa_s0_c22_n43_s),
        .c_out(fa_s0_c22_n43_c)
    );

    fa fa_s0_c23_n44 (
        .a(stage0_col23[0]),
        .b(stage0_col23[1]),
        .c_in(stage0_col23[2]),
        .s(fa_s0_c23_n44_s),
        .c_out(fa_s0_c23_n44_c)
    );

    fa fa_s0_c23_n45 (
        .a(stage0_col23[3]),
        .b(stage0_col23[4]),
        .c_in(stage0_col23[5]),
        .s(fa_s0_c23_n45_s),
        .c_out(fa_s0_c23_n45_c)
    );

    fa fa_s0_c23_n46 (
        .a(stage0_col23[6]),
        .b(stage0_col23[7]),
        .c_in(stage0_col23[8]),
        .s(fa_s0_c23_n46_s),
        .c_out(fa_s0_c23_n46_c)
    );

    fa fa_s0_c23_n47 (
        .a(stage0_col23[9]),
        .b(stage0_col23[10]),
        .c_in(stage0_col23[11]),
        .s(fa_s0_c23_n47_s),
        .c_out(fa_s0_c23_n47_c)
    );

    fa fa_s0_c24_n48 (
        .a(stage0_col24[0]),
        .b(stage0_col24[1]),
        .c_in(stage0_col24[2]),
        .s(fa_s0_c24_n48_s),
        .c_out(fa_s0_c24_n48_c)
    );

    fa fa_s0_c24_n49 (
        .a(stage0_col24[3]),
        .b(stage0_col24[4]),
        .c_in(stage0_col24[5]),
        .s(fa_s0_c24_n49_s),
        .c_out(fa_s0_c24_n49_c)
    );

    fa fa_s0_c24_n50 (
        .a(stage0_col24[6]),
        .b(stage0_col24[7]),
        .c_in(stage0_col24[8]),
        .s(fa_s0_c24_n50_s),
        .c_out(fa_s0_c24_n50_c)
    );

    fa fa_s0_c24_n51 (
        .a(stage0_col24[9]),
        .b(stage0_col24[10]),
        .c_in(stage0_col24[11]),
        .s(fa_s0_c24_n51_s),
        .c_out(fa_s0_c24_n51_c)
    );

    fa fa_s0_c25_n52 (
        .a(stage0_col25[0]),
        .b(stage0_col25[1]),
        .c_in(stage0_col25[2]),
        .s(fa_s0_c25_n52_s),
        .c_out(fa_s0_c25_n52_c)
    );

    fa fa_s0_c25_n53 (
        .a(stage0_col25[3]),
        .b(stage0_col25[4]),
        .c_in(stage0_col25[5]),
        .s(fa_s0_c25_n53_s),
        .c_out(fa_s0_c25_n53_c)
    );

    fa fa_s0_c25_n54 (
        .a(stage0_col25[6]),
        .b(stage0_col25[7]),
        .c_in(stage0_col25[8]),
        .s(fa_s0_c25_n54_s),
        .c_out(fa_s0_c25_n54_c)
    );

    fa fa_s0_c25_n55 (
        .a(stage0_col25[9]),
        .b(stage0_col25[10]),
        .c_in(stage0_col25[11]),
        .s(fa_s0_c25_n55_s),
        .c_out(fa_s0_c25_n55_c)
    );

    fa fa_s0_c26_n56 (
        .a(stage0_col26[0]),
        .b(stage0_col26[1]),
        .c_in(stage0_col26[2]),
        .s(fa_s0_c26_n56_s),
        .c_out(fa_s0_c26_n56_c)
    );

    fa fa_s0_c26_n57 (
        .a(stage0_col26[3]),
        .b(stage0_col26[4]),
        .c_in(stage0_col26[5]),
        .s(fa_s0_c26_n57_s),
        .c_out(fa_s0_c26_n57_c)
    );

    fa fa_s0_c26_n58 (
        .a(stage0_col26[6]),
        .b(stage0_col26[7]),
        .c_in(stage0_col26[8]),
        .s(fa_s0_c26_n58_s),
        .c_out(fa_s0_c26_n58_c)
    );

    fa fa_s0_c26_n59 (
        .a(stage0_col26[9]),
        .b(stage0_col26[10]),
        .c_in(stage0_col26[11]),
        .s(fa_s0_c26_n59_s),
        .c_out(fa_s0_c26_n59_c)
    );

    fa fa_s0_c26_n60 (
        .a(stage0_col26[12]),
        .b(stage0_col26[13]),
        .c_in(stage0_col26[14]),
        .s(fa_s0_c26_n60_s),
        .c_out(fa_s0_c26_n60_c)
    );

    fa fa_s0_c27_n61 (
        .a(stage0_col27[0]),
        .b(stage0_col27[1]),
        .c_in(stage0_col27[2]),
        .s(fa_s0_c27_n61_s),
        .c_out(fa_s0_c27_n61_c)
    );

    fa fa_s0_c27_n62 (
        .a(stage0_col27[3]),
        .b(stage0_col27[4]),
        .c_in(stage0_col27[5]),
        .s(fa_s0_c27_n62_s),
        .c_out(fa_s0_c27_n62_c)
    );

    fa fa_s0_c27_n63 (
        .a(stage0_col27[6]),
        .b(stage0_col27[7]),
        .c_in(stage0_col27[8]),
        .s(fa_s0_c27_n63_s),
        .c_out(fa_s0_c27_n63_c)
    );

    fa fa_s0_c27_n64 (
        .a(stage0_col27[9]),
        .b(stage0_col27[10]),
        .c_in(stage0_col27[11]),
        .s(fa_s0_c27_n64_s),
        .c_out(fa_s0_c27_n64_c)
    );

    fa fa_s0_c28_n65 (
        .a(stage0_col28[0]),
        .b(stage0_col28[1]),
        .c_in(stage0_col28[2]),
        .s(fa_s0_c28_n65_s),
        .c_out(fa_s0_c28_n65_c)
    );

    fa fa_s0_c28_n66 (
        .a(stage0_col28[3]),
        .b(stage0_col28[4]),
        .c_in(stage0_col28[5]),
        .s(fa_s0_c28_n66_s),
        .c_out(fa_s0_c28_n66_c)
    );

    fa fa_s0_c28_n67 (
        .a(stage0_col28[6]),
        .b(stage0_col28[7]),
        .c_in(stage0_col28[8]),
        .s(fa_s0_c28_n67_s),
        .c_out(fa_s0_c28_n67_c)
    );

    fa fa_s0_c28_n68 (
        .a(stage0_col28[9]),
        .b(stage0_col28[10]),
        .c_in(stage0_col28[11]),
        .s(fa_s0_c28_n68_s),
        .c_out(fa_s0_c28_n68_c)
    );

    fa fa_s0_c28_n69 (
        .a(stage0_col28[12]),
        .b(stage0_col28[13]),
        .c_in(stage0_col28[14]),
        .s(fa_s0_c28_n69_s),
        .c_out(fa_s0_c28_n69_c)
    );

    fa fa_s0_c29_n70 (
        .a(stage0_col29[0]),
        .b(stage0_col29[1]),
        .c_in(stage0_col29[2]),
        .s(fa_s0_c29_n70_s),
        .c_out(fa_s0_c29_n70_c)
    );

    fa fa_s0_c29_n71 (
        .a(stage0_col29[3]),
        .b(stage0_col29[4]),
        .c_in(stage0_col29[5]),
        .s(fa_s0_c29_n71_s),
        .c_out(fa_s0_c29_n71_c)
    );

    fa fa_s0_c29_n72 (
        .a(stage0_col29[6]),
        .b(stage0_col29[7]),
        .c_in(stage0_col29[8]),
        .s(fa_s0_c29_n72_s),
        .c_out(fa_s0_c29_n72_c)
    );

    fa fa_s0_c29_n73 (
        .a(stage0_col29[9]),
        .b(stage0_col29[10]),
        .c_in(stage0_col29[11]),
        .s(fa_s0_c29_n73_s),
        .c_out(fa_s0_c29_n73_c)
    );

    fa fa_s0_c29_n74 (
        .a(stage0_col29[12]),
        .b(stage0_col29[13]),
        .c_in(stage0_col29[14]),
        .s(fa_s0_c29_n74_s),
        .c_out(fa_s0_c29_n74_c)
    );

    fa fa_s0_c30_n75 (
        .a(stage0_col30[0]),
        .b(stage0_col30[1]),
        .c_in(stage0_col30[2]),
        .s(fa_s0_c30_n75_s),
        .c_out(fa_s0_c30_n75_c)
    );

    fa fa_s0_c30_n76 (
        .a(stage0_col30[3]),
        .b(stage0_col30[4]),
        .c_in(stage0_col30[5]),
        .s(fa_s0_c30_n76_s),
        .c_out(fa_s0_c30_n76_c)
    );

    fa fa_s0_c30_n77 (
        .a(stage0_col30[6]),
        .b(stage0_col30[7]),
        .c_in(stage0_col30[8]),
        .s(fa_s0_c30_n77_s),
        .c_out(fa_s0_c30_n77_c)
    );

    fa fa_s0_c30_n78 (
        .a(stage0_col30[9]),
        .b(stage0_col30[10]),
        .c_in(stage0_col30[11]),
        .s(fa_s0_c30_n78_s),
        .c_out(fa_s0_c30_n78_c)
    );

    fa fa_s0_c30_n79 (
        .a(stage0_col30[12]),
        .b(stage0_col30[13]),
        .c_in(stage0_col30[14]),
        .s(fa_s0_c30_n79_s),
        .c_out(fa_s0_c30_n79_c)
    );

    fa fa_s0_c31_n80 (
        .a(stage0_col31[0]),
        .b(stage0_col31[1]),
        .c_in(stage0_col31[2]),
        .s(fa_s0_c31_n80_s),
        .c_out(fa_s0_c31_n80_c)
    );

    fa fa_s0_c31_n81 (
        .a(stage0_col31[3]),
        .b(stage0_col31[4]),
        .c_in(stage0_col31[5]),
        .s(fa_s0_c31_n81_s),
        .c_out(fa_s0_c31_n81_c)
    );

    fa fa_s0_c31_n82 (
        .a(stage0_col31[6]),
        .b(stage0_col31[7]),
        .c_in(stage0_col31[8]),
        .s(fa_s0_c31_n82_s),
        .c_out(fa_s0_c31_n82_c)
    );

    fa fa_s0_c31_n83 (
        .a(stage0_col31[9]),
        .b(stage0_col31[10]),
        .c_in(stage0_col31[11]),
        .s(fa_s0_c31_n83_s),
        .c_out(fa_s0_c31_n83_c)
    );

    fa fa_s0_c31_n84 (
        .a(stage0_col31[12]),
        .b(stage0_col31[13]),
        .c_in(stage0_col31[14]),
        .s(fa_s0_c31_n84_s),
        .c_out(fa_s0_c31_n84_c)
    );

    fa fa_s0_c32_n85 (
        .a(stage0_col32[0]),
        .b(stage0_col32[1]),
        .c_in(stage0_col32[2]),
        .s(fa_s0_c32_n85_s),
        .c_out(fa_s0_c32_n85_c)
    );

    fa fa_s0_c32_n86 (
        .a(stage0_col32[3]),
        .b(stage0_col32[4]),
        .c_in(stage0_col32[5]),
        .s(fa_s0_c32_n86_s),
        .c_out(fa_s0_c32_n86_c)
    );

    fa fa_s0_c32_n87 (
        .a(stage0_col32[6]),
        .b(stage0_col32[7]),
        .c_in(stage0_col32[8]),
        .s(fa_s0_c32_n87_s),
        .c_out(fa_s0_c32_n87_c)
    );

    fa fa_s0_c32_n88 (
        .a(stage0_col32[9]),
        .b(stage0_col32[10]),
        .c_in(stage0_col32[11]),
        .s(fa_s0_c32_n88_s),
        .c_out(fa_s0_c32_n88_c)
    );

    fa fa_s0_c32_n89 (
        .a(stage0_col32[12]),
        .b(stage0_col32[13]),
        .c_in(stage0_col32[14]),
        .s(fa_s0_c32_n89_s),
        .c_out(fa_s0_c32_n89_c)
    );

    fa fa_s0_c32_n90 (
        .a(stage0_col32[15]),
        .b(stage0_col32[16]),
        .c_in(stage0_col32[17]),
        .s(fa_s0_c32_n90_s),
        .c_out(fa_s0_c32_n90_c)
    );

    fa fa_s0_c33_n91 (
        .a(stage0_col33[0]),
        .b(stage0_col33[1]),
        .c_in(stage0_col33[2]),
        .s(fa_s0_c33_n91_s),
        .c_out(fa_s0_c33_n91_c)
    );

    fa fa_s0_c33_n92 (
        .a(stage0_col33[3]),
        .b(stage0_col33[4]),
        .c_in(stage0_col33[5]),
        .s(fa_s0_c33_n92_s),
        .c_out(fa_s0_c33_n92_c)
    );

    fa fa_s0_c33_n93 (
        .a(stage0_col33[6]),
        .b(stage0_col33[7]),
        .c_in(stage0_col33[8]),
        .s(fa_s0_c33_n93_s),
        .c_out(fa_s0_c33_n93_c)
    );

    fa fa_s0_c33_n94 (
        .a(stage0_col33[9]),
        .b(stage0_col33[10]),
        .c_in(stage0_col33[11]),
        .s(fa_s0_c33_n94_s),
        .c_out(fa_s0_c33_n94_c)
    );

    fa fa_s0_c33_n95 (
        .a(stage0_col33[12]),
        .b(stage0_col33[13]),
        .c_in(stage0_col33[14]),
        .s(fa_s0_c33_n95_s),
        .c_out(fa_s0_c33_n95_c)
    );

    fa fa_s0_c34_n96 (
        .a(stage0_col34[0]),
        .b(stage0_col34[1]),
        .c_in(stage0_col34[2]),
        .s(fa_s0_c34_n96_s),
        .c_out(fa_s0_c34_n96_c)
    );

    fa fa_s0_c34_n97 (
        .a(stage0_col34[3]),
        .b(stage0_col34[4]),
        .c_in(stage0_col34[5]),
        .s(fa_s0_c34_n97_s),
        .c_out(fa_s0_c34_n97_c)
    );

    fa fa_s0_c34_n98 (
        .a(stage0_col34[6]),
        .b(stage0_col34[7]),
        .c_in(stage0_col34[8]),
        .s(fa_s0_c34_n98_s),
        .c_out(fa_s0_c34_n98_c)
    );

    fa fa_s0_c34_n99 (
        .a(stage0_col34[9]),
        .b(stage0_col34[10]),
        .c_in(stage0_col34[11]),
        .s(fa_s0_c34_n99_s),
        .c_out(fa_s0_c34_n99_c)
    );

    fa fa_s0_c34_n100 (
        .a(stage0_col34[12]),
        .b(stage0_col34[13]),
        .c_in(stage0_col34[14]),
        .s(fa_s0_c34_n100_s),
        .c_out(fa_s0_c34_n100_c)
    );

    fa fa_s0_c34_n101 (
        .a(stage0_col34[15]),
        .b(stage0_col34[16]),
        .c_in(stage0_col34[17]),
        .s(fa_s0_c34_n101_s),
        .c_out(fa_s0_c34_n101_c)
    );

    fa fa_s0_c35_n102 (
        .a(stage0_col35[0]),
        .b(stage0_col35[1]),
        .c_in(stage0_col35[2]),
        .s(fa_s0_c35_n102_s),
        .c_out(fa_s0_c35_n102_c)
    );

    fa fa_s0_c35_n103 (
        .a(stage0_col35[3]),
        .b(stage0_col35[4]),
        .c_in(stage0_col35[5]),
        .s(fa_s0_c35_n103_s),
        .c_out(fa_s0_c35_n103_c)
    );

    fa fa_s0_c35_n104 (
        .a(stage0_col35[6]),
        .b(stage0_col35[7]),
        .c_in(stage0_col35[8]),
        .s(fa_s0_c35_n104_s),
        .c_out(fa_s0_c35_n104_c)
    );

    fa fa_s0_c35_n105 (
        .a(stage0_col35[9]),
        .b(stage0_col35[10]),
        .c_in(stage0_col35[11]),
        .s(fa_s0_c35_n105_s),
        .c_out(fa_s0_c35_n105_c)
    );

    fa fa_s0_c35_n106 (
        .a(stage0_col35[12]),
        .b(stage0_col35[13]),
        .c_in(stage0_col35[14]),
        .s(fa_s0_c35_n106_s),
        .c_out(fa_s0_c35_n106_c)
    );

    fa fa_s0_c35_n107 (
        .a(stage0_col35[15]),
        .b(stage0_col35[16]),
        .c_in(stage0_col35[17]),
        .s(fa_s0_c35_n107_s),
        .c_out(fa_s0_c35_n107_c)
    );

    fa fa_s0_c36_n108 (
        .a(stage0_col36[0]),
        .b(stage0_col36[1]),
        .c_in(stage0_col36[2]),
        .s(fa_s0_c36_n108_s),
        .c_out(fa_s0_c36_n108_c)
    );

    fa fa_s0_c36_n109 (
        .a(stage0_col36[3]),
        .b(stage0_col36[4]),
        .c_in(stage0_col36[5]),
        .s(fa_s0_c36_n109_s),
        .c_out(fa_s0_c36_n109_c)
    );

    fa fa_s0_c36_n110 (
        .a(stage0_col36[6]),
        .b(stage0_col36[7]),
        .c_in(stage0_col36[8]),
        .s(fa_s0_c36_n110_s),
        .c_out(fa_s0_c36_n110_c)
    );

    fa fa_s0_c36_n111 (
        .a(stage0_col36[9]),
        .b(stage0_col36[10]),
        .c_in(stage0_col36[11]),
        .s(fa_s0_c36_n111_s),
        .c_out(fa_s0_c36_n111_c)
    );

    fa fa_s0_c36_n112 (
        .a(stage0_col36[12]),
        .b(stage0_col36[13]),
        .c_in(stage0_col36[14]),
        .s(fa_s0_c36_n112_s),
        .c_out(fa_s0_c36_n112_c)
    );

    fa fa_s0_c36_n113 (
        .a(stage0_col36[15]),
        .b(stage0_col36[16]),
        .c_in(stage0_col36[17]),
        .s(fa_s0_c36_n113_s),
        .c_out(fa_s0_c36_n113_c)
    );

    fa fa_s0_c37_n114 (
        .a(stage0_col37[0]),
        .b(stage0_col37[1]),
        .c_in(stage0_col37[2]),
        .s(fa_s0_c37_n114_s),
        .c_out(fa_s0_c37_n114_c)
    );

    fa fa_s0_c37_n115 (
        .a(stage0_col37[3]),
        .b(stage0_col37[4]),
        .c_in(stage0_col37[5]),
        .s(fa_s0_c37_n115_s),
        .c_out(fa_s0_c37_n115_c)
    );

    fa fa_s0_c37_n116 (
        .a(stage0_col37[6]),
        .b(stage0_col37[7]),
        .c_in(stage0_col37[8]),
        .s(fa_s0_c37_n116_s),
        .c_out(fa_s0_c37_n116_c)
    );

    fa fa_s0_c37_n117 (
        .a(stage0_col37[9]),
        .b(stage0_col37[10]),
        .c_in(stage0_col37[11]),
        .s(fa_s0_c37_n117_s),
        .c_out(fa_s0_c37_n117_c)
    );

    fa fa_s0_c37_n118 (
        .a(stage0_col37[12]),
        .b(stage0_col37[13]),
        .c_in(stage0_col37[14]),
        .s(fa_s0_c37_n118_s),
        .c_out(fa_s0_c37_n118_c)
    );

    fa fa_s0_c37_n119 (
        .a(stage0_col37[15]),
        .b(stage0_col37[16]),
        .c_in(stage0_col37[17]),
        .s(fa_s0_c37_n119_s),
        .c_out(fa_s0_c37_n119_c)
    );

    fa fa_s0_c38_n120 (
        .a(stage0_col38[0]),
        .b(stage0_col38[1]),
        .c_in(stage0_col38[2]),
        .s(fa_s0_c38_n120_s),
        .c_out(fa_s0_c38_n120_c)
    );

    fa fa_s0_c38_n121 (
        .a(stage0_col38[3]),
        .b(stage0_col38[4]),
        .c_in(stage0_col38[5]),
        .s(fa_s0_c38_n121_s),
        .c_out(fa_s0_c38_n121_c)
    );

    fa fa_s0_c38_n122 (
        .a(stage0_col38[6]),
        .b(stage0_col38[7]),
        .c_in(stage0_col38[8]),
        .s(fa_s0_c38_n122_s),
        .c_out(fa_s0_c38_n122_c)
    );

    fa fa_s0_c38_n123 (
        .a(stage0_col38[9]),
        .b(stage0_col38[10]),
        .c_in(stage0_col38[11]),
        .s(fa_s0_c38_n123_s),
        .c_out(fa_s0_c38_n123_c)
    );

    fa fa_s0_c38_n124 (
        .a(stage0_col38[12]),
        .b(stage0_col38[13]),
        .c_in(stage0_col38[14]),
        .s(fa_s0_c38_n124_s),
        .c_out(fa_s0_c38_n124_c)
    );

    fa fa_s0_c38_n125 (
        .a(stage0_col38[15]),
        .b(stage0_col38[16]),
        .c_in(stage0_col38[17]),
        .s(fa_s0_c38_n125_s),
        .c_out(fa_s0_c38_n125_c)
    );

    fa fa_s0_c38_n126 (
        .a(stage0_col38[18]),
        .b(stage0_col38[19]),
        .c_in(stage0_col38[20]),
        .s(fa_s0_c38_n126_s),
        .c_out(fa_s0_c38_n126_c)
    );

    fa fa_s0_c39_n127 (
        .a(stage0_col39[0]),
        .b(stage0_col39[1]),
        .c_in(stage0_col39[2]),
        .s(fa_s0_c39_n127_s),
        .c_out(fa_s0_c39_n127_c)
    );

    fa fa_s0_c39_n128 (
        .a(stage0_col39[3]),
        .b(stage0_col39[4]),
        .c_in(stage0_col39[5]),
        .s(fa_s0_c39_n128_s),
        .c_out(fa_s0_c39_n128_c)
    );

    fa fa_s0_c39_n129 (
        .a(stage0_col39[6]),
        .b(stage0_col39[7]),
        .c_in(stage0_col39[8]),
        .s(fa_s0_c39_n129_s),
        .c_out(fa_s0_c39_n129_c)
    );

    fa fa_s0_c39_n130 (
        .a(stage0_col39[9]),
        .b(stage0_col39[10]),
        .c_in(stage0_col39[11]),
        .s(fa_s0_c39_n130_s),
        .c_out(fa_s0_c39_n130_c)
    );

    fa fa_s0_c39_n131 (
        .a(stage0_col39[12]),
        .b(stage0_col39[13]),
        .c_in(stage0_col39[14]),
        .s(fa_s0_c39_n131_s),
        .c_out(fa_s0_c39_n131_c)
    );

    fa fa_s0_c39_n132 (
        .a(stage0_col39[15]),
        .b(stage0_col39[16]),
        .c_in(stage0_col39[17]),
        .s(fa_s0_c39_n132_s),
        .c_out(fa_s0_c39_n132_c)
    );

    fa fa_s0_c40_n133 (
        .a(stage0_col40[0]),
        .b(stage0_col40[1]),
        .c_in(stage0_col40[2]),
        .s(fa_s0_c40_n133_s),
        .c_out(fa_s0_c40_n133_c)
    );

    fa fa_s0_c40_n134 (
        .a(stage0_col40[3]),
        .b(stage0_col40[4]),
        .c_in(stage0_col40[5]),
        .s(fa_s0_c40_n134_s),
        .c_out(fa_s0_c40_n134_c)
    );

    fa fa_s0_c40_n135 (
        .a(stage0_col40[6]),
        .b(stage0_col40[7]),
        .c_in(stage0_col40[8]),
        .s(fa_s0_c40_n135_s),
        .c_out(fa_s0_c40_n135_c)
    );

    fa fa_s0_c40_n136 (
        .a(stage0_col40[9]),
        .b(stage0_col40[10]),
        .c_in(stage0_col40[11]),
        .s(fa_s0_c40_n136_s),
        .c_out(fa_s0_c40_n136_c)
    );

    fa fa_s0_c40_n137 (
        .a(stage0_col40[12]),
        .b(stage0_col40[13]),
        .c_in(stage0_col40[14]),
        .s(fa_s0_c40_n137_s),
        .c_out(fa_s0_c40_n137_c)
    );

    fa fa_s0_c40_n138 (
        .a(stage0_col40[15]),
        .b(stage0_col40[16]),
        .c_in(stage0_col40[17]),
        .s(fa_s0_c40_n138_s),
        .c_out(fa_s0_c40_n138_c)
    );

    fa fa_s0_c40_n139 (
        .a(stage0_col40[18]),
        .b(stage0_col40[19]),
        .c_in(stage0_col40[20]),
        .s(fa_s0_c40_n139_s),
        .c_out(fa_s0_c40_n139_c)
    );

    fa fa_s0_c41_n140 (
        .a(stage0_col41[0]),
        .b(stage0_col41[1]),
        .c_in(stage0_col41[2]),
        .s(fa_s0_c41_n140_s),
        .c_out(fa_s0_c41_n140_c)
    );

    fa fa_s0_c41_n141 (
        .a(stage0_col41[3]),
        .b(stage0_col41[4]),
        .c_in(stage0_col41[5]),
        .s(fa_s0_c41_n141_s),
        .c_out(fa_s0_c41_n141_c)
    );

    fa fa_s0_c41_n142 (
        .a(stage0_col41[6]),
        .b(stage0_col41[7]),
        .c_in(stage0_col41[8]),
        .s(fa_s0_c41_n142_s),
        .c_out(fa_s0_c41_n142_c)
    );

    fa fa_s0_c41_n143 (
        .a(stage0_col41[9]),
        .b(stage0_col41[10]),
        .c_in(stage0_col41[11]),
        .s(fa_s0_c41_n143_s),
        .c_out(fa_s0_c41_n143_c)
    );

    fa fa_s0_c41_n144 (
        .a(stage0_col41[12]),
        .b(stage0_col41[13]),
        .c_in(stage0_col41[14]),
        .s(fa_s0_c41_n144_s),
        .c_out(fa_s0_c41_n144_c)
    );

    fa fa_s0_c41_n145 (
        .a(stage0_col41[15]),
        .b(stage0_col41[16]),
        .c_in(stage0_col41[17]),
        .s(fa_s0_c41_n145_s),
        .c_out(fa_s0_c41_n145_c)
    );

    fa fa_s0_c41_n146 (
        .a(stage0_col41[18]),
        .b(stage0_col41[19]),
        .c_in(stage0_col41[20]),
        .s(fa_s0_c41_n146_s),
        .c_out(fa_s0_c41_n146_c)
    );

    fa fa_s0_c42_n147 (
        .a(stage0_col42[0]),
        .b(stage0_col42[1]),
        .c_in(stage0_col42[2]),
        .s(fa_s0_c42_n147_s),
        .c_out(fa_s0_c42_n147_c)
    );

    fa fa_s0_c42_n148 (
        .a(stage0_col42[3]),
        .b(stage0_col42[4]),
        .c_in(stage0_col42[5]),
        .s(fa_s0_c42_n148_s),
        .c_out(fa_s0_c42_n148_c)
    );

    fa fa_s0_c42_n149 (
        .a(stage0_col42[6]),
        .b(stage0_col42[7]),
        .c_in(stage0_col42[8]),
        .s(fa_s0_c42_n149_s),
        .c_out(fa_s0_c42_n149_c)
    );

    fa fa_s0_c42_n150 (
        .a(stage0_col42[9]),
        .b(stage0_col42[10]),
        .c_in(stage0_col42[11]),
        .s(fa_s0_c42_n150_s),
        .c_out(fa_s0_c42_n150_c)
    );

    fa fa_s0_c42_n151 (
        .a(stage0_col42[12]),
        .b(stage0_col42[13]),
        .c_in(stage0_col42[14]),
        .s(fa_s0_c42_n151_s),
        .c_out(fa_s0_c42_n151_c)
    );

    fa fa_s0_c42_n152 (
        .a(stage0_col42[15]),
        .b(stage0_col42[16]),
        .c_in(stage0_col42[17]),
        .s(fa_s0_c42_n152_s),
        .c_out(fa_s0_c42_n152_c)
    );

    fa fa_s0_c42_n153 (
        .a(stage0_col42[18]),
        .b(stage0_col42[19]),
        .c_in(stage0_col42[20]),
        .s(fa_s0_c42_n153_s),
        .c_out(fa_s0_c42_n153_c)
    );

    fa fa_s0_c43_n154 (
        .a(stage0_col43[0]),
        .b(stage0_col43[1]),
        .c_in(stage0_col43[2]),
        .s(fa_s0_c43_n154_s),
        .c_out(fa_s0_c43_n154_c)
    );

    fa fa_s0_c43_n155 (
        .a(stage0_col43[3]),
        .b(stage0_col43[4]),
        .c_in(stage0_col43[5]),
        .s(fa_s0_c43_n155_s),
        .c_out(fa_s0_c43_n155_c)
    );

    fa fa_s0_c43_n156 (
        .a(stage0_col43[6]),
        .b(stage0_col43[7]),
        .c_in(stage0_col43[8]),
        .s(fa_s0_c43_n156_s),
        .c_out(fa_s0_c43_n156_c)
    );

    fa fa_s0_c43_n157 (
        .a(stage0_col43[9]),
        .b(stage0_col43[10]),
        .c_in(stage0_col43[11]),
        .s(fa_s0_c43_n157_s),
        .c_out(fa_s0_c43_n157_c)
    );

    fa fa_s0_c43_n158 (
        .a(stage0_col43[12]),
        .b(stage0_col43[13]),
        .c_in(stage0_col43[14]),
        .s(fa_s0_c43_n158_s),
        .c_out(fa_s0_c43_n158_c)
    );

    fa fa_s0_c43_n159 (
        .a(stage0_col43[15]),
        .b(stage0_col43[16]),
        .c_in(stage0_col43[17]),
        .s(fa_s0_c43_n159_s),
        .c_out(fa_s0_c43_n159_c)
    );

    fa fa_s0_c43_n160 (
        .a(stage0_col43[18]),
        .b(stage0_col43[19]),
        .c_in(stage0_col43[20]),
        .s(fa_s0_c43_n160_s),
        .c_out(fa_s0_c43_n160_c)
    );

    fa fa_s0_c44_n161 (
        .a(stage0_col44[0]),
        .b(stage0_col44[1]),
        .c_in(stage0_col44[2]),
        .s(fa_s0_c44_n161_s),
        .c_out(fa_s0_c44_n161_c)
    );

    fa fa_s0_c44_n162 (
        .a(stage0_col44[3]),
        .b(stage0_col44[4]),
        .c_in(stage0_col44[5]),
        .s(fa_s0_c44_n162_s),
        .c_out(fa_s0_c44_n162_c)
    );

    fa fa_s0_c44_n163 (
        .a(stage0_col44[6]),
        .b(stage0_col44[7]),
        .c_in(stage0_col44[8]),
        .s(fa_s0_c44_n163_s),
        .c_out(fa_s0_c44_n163_c)
    );

    fa fa_s0_c44_n164 (
        .a(stage0_col44[9]),
        .b(stage0_col44[10]),
        .c_in(stage0_col44[11]),
        .s(fa_s0_c44_n164_s),
        .c_out(fa_s0_c44_n164_c)
    );

    fa fa_s0_c44_n165 (
        .a(stage0_col44[12]),
        .b(stage0_col44[13]),
        .c_in(stage0_col44[14]),
        .s(fa_s0_c44_n165_s),
        .c_out(fa_s0_c44_n165_c)
    );

    fa fa_s0_c44_n166 (
        .a(stage0_col44[15]),
        .b(stage0_col44[16]),
        .c_in(stage0_col44[17]),
        .s(fa_s0_c44_n166_s),
        .c_out(fa_s0_c44_n166_c)
    );

    fa fa_s0_c44_n167 (
        .a(stage0_col44[18]),
        .b(stage0_col44[19]),
        .c_in(stage0_col44[20]),
        .s(fa_s0_c44_n167_s),
        .c_out(fa_s0_c44_n167_c)
    );

    fa fa_s0_c44_n168 (
        .a(stage0_col44[21]),
        .b(stage0_col44[22]),
        .c_in(stage0_col44[23]),
        .s(fa_s0_c44_n168_s),
        .c_out(fa_s0_c44_n168_c)
    );

    fa fa_s0_c45_n169 (
        .a(stage0_col45[0]),
        .b(stage0_col45[1]),
        .c_in(stage0_col45[2]),
        .s(fa_s0_c45_n169_s),
        .c_out(fa_s0_c45_n169_c)
    );

    fa fa_s0_c45_n170 (
        .a(stage0_col45[3]),
        .b(stage0_col45[4]),
        .c_in(stage0_col45[5]),
        .s(fa_s0_c45_n170_s),
        .c_out(fa_s0_c45_n170_c)
    );

    fa fa_s0_c45_n171 (
        .a(stage0_col45[6]),
        .b(stage0_col45[7]),
        .c_in(stage0_col45[8]),
        .s(fa_s0_c45_n171_s),
        .c_out(fa_s0_c45_n171_c)
    );

    fa fa_s0_c45_n172 (
        .a(stage0_col45[9]),
        .b(stage0_col45[10]),
        .c_in(stage0_col45[11]),
        .s(fa_s0_c45_n172_s),
        .c_out(fa_s0_c45_n172_c)
    );

    fa fa_s0_c45_n173 (
        .a(stage0_col45[12]),
        .b(stage0_col45[13]),
        .c_in(stage0_col45[14]),
        .s(fa_s0_c45_n173_s),
        .c_out(fa_s0_c45_n173_c)
    );

    fa fa_s0_c45_n174 (
        .a(stage0_col45[15]),
        .b(stage0_col45[16]),
        .c_in(stage0_col45[17]),
        .s(fa_s0_c45_n174_s),
        .c_out(fa_s0_c45_n174_c)
    );

    fa fa_s0_c45_n175 (
        .a(stage0_col45[18]),
        .b(stage0_col45[19]),
        .c_in(stage0_col45[20]),
        .s(fa_s0_c45_n175_s),
        .c_out(fa_s0_c45_n175_c)
    );

    fa fa_s0_c46_n176 (
        .a(stage0_col46[0]),
        .b(stage0_col46[1]),
        .c_in(stage0_col46[2]),
        .s(fa_s0_c46_n176_s),
        .c_out(fa_s0_c46_n176_c)
    );

    fa fa_s0_c46_n177 (
        .a(stage0_col46[3]),
        .b(stage0_col46[4]),
        .c_in(stage0_col46[5]),
        .s(fa_s0_c46_n177_s),
        .c_out(fa_s0_c46_n177_c)
    );

    fa fa_s0_c46_n178 (
        .a(stage0_col46[6]),
        .b(stage0_col46[7]),
        .c_in(stage0_col46[8]),
        .s(fa_s0_c46_n178_s),
        .c_out(fa_s0_c46_n178_c)
    );

    fa fa_s0_c46_n179 (
        .a(stage0_col46[9]),
        .b(stage0_col46[10]),
        .c_in(stage0_col46[11]),
        .s(fa_s0_c46_n179_s),
        .c_out(fa_s0_c46_n179_c)
    );

    fa fa_s0_c46_n180 (
        .a(stage0_col46[12]),
        .b(stage0_col46[13]),
        .c_in(stage0_col46[14]),
        .s(fa_s0_c46_n180_s),
        .c_out(fa_s0_c46_n180_c)
    );

    fa fa_s0_c46_n181 (
        .a(stage0_col46[15]),
        .b(stage0_col46[16]),
        .c_in(stage0_col46[17]),
        .s(fa_s0_c46_n181_s),
        .c_out(fa_s0_c46_n181_c)
    );

    fa fa_s0_c46_n182 (
        .a(stage0_col46[18]),
        .b(stage0_col46[19]),
        .c_in(stage0_col46[20]),
        .s(fa_s0_c46_n182_s),
        .c_out(fa_s0_c46_n182_c)
    );

    fa fa_s0_c46_n183 (
        .a(stage0_col46[21]),
        .b(stage0_col46[22]),
        .c_in(stage0_col46[23]),
        .s(fa_s0_c46_n183_s),
        .c_out(fa_s0_c46_n183_c)
    );

    fa fa_s0_c47_n184 (
        .a(stage0_col47[0]),
        .b(stage0_col47[1]),
        .c_in(stage0_col47[2]),
        .s(fa_s0_c47_n184_s),
        .c_out(fa_s0_c47_n184_c)
    );

    fa fa_s0_c47_n185 (
        .a(stage0_col47[3]),
        .b(stage0_col47[4]),
        .c_in(stage0_col47[5]),
        .s(fa_s0_c47_n185_s),
        .c_out(fa_s0_c47_n185_c)
    );

    fa fa_s0_c47_n186 (
        .a(stage0_col47[6]),
        .b(stage0_col47[7]),
        .c_in(stage0_col47[8]),
        .s(fa_s0_c47_n186_s),
        .c_out(fa_s0_c47_n186_c)
    );

    fa fa_s0_c47_n187 (
        .a(stage0_col47[9]),
        .b(stage0_col47[10]),
        .c_in(stage0_col47[11]),
        .s(fa_s0_c47_n187_s),
        .c_out(fa_s0_c47_n187_c)
    );

    fa fa_s0_c47_n188 (
        .a(stage0_col47[12]),
        .b(stage0_col47[13]),
        .c_in(stage0_col47[14]),
        .s(fa_s0_c47_n188_s),
        .c_out(fa_s0_c47_n188_c)
    );

    fa fa_s0_c47_n189 (
        .a(stage0_col47[15]),
        .b(stage0_col47[16]),
        .c_in(stage0_col47[17]),
        .s(fa_s0_c47_n189_s),
        .c_out(fa_s0_c47_n189_c)
    );

    fa fa_s0_c47_n190 (
        .a(stage0_col47[18]),
        .b(stage0_col47[19]),
        .c_in(stage0_col47[20]),
        .s(fa_s0_c47_n190_s),
        .c_out(fa_s0_c47_n190_c)
    );

    fa fa_s0_c47_n191 (
        .a(stage0_col47[21]),
        .b(stage0_col47[22]),
        .c_in(stage0_col47[23]),
        .s(fa_s0_c47_n191_s),
        .c_out(fa_s0_c47_n191_c)
    );

    fa fa_s0_c48_n192 (
        .a(stage0_col48[0]),
        .b(stage0_col48[1]),
        .c_in(stage0_col48[2]),
        .s(fa_s0_c48_n192_s),
        .c_out(fa_s0_c48_n192_c)
    );

    fa fa_s0_c48_n193 (
        .a(stage0_col48[3]),
        .b(stage0_col48[4]),
        .c_in(stage0_col48[5]),
        .s(fa_s0_c48_n193_s),
        .c_out(fa_s0_c48_n193_c)
    );

    fa fa_s0_c48_n194 (
        .a(stage0_col48[6]),
        .b(stage0_col48[7]),
        .c_in(stage0_col48[8]),
        .s(fa_s0_c48_n194_s),
        .c_out(fa_s0_c48_n194_c)
    );

    fa fa_s0_c48_n195 (
        .a(stage0_col48[9]),
        .b(stage0_col48[10]),
        .c_in(stage0_col48[11]),
        .s(fa_s0_c48_n195_s),
        .c_out(fa_s0_c48_n195_c)
    );

    fa fa_s0_c48_n196 (
        .a(stage0_col48[12]),
        .b(stage0_col48[13]),
        .c_in(stage0_col48[14]),
        .s(fa_s0_c48_n196_s),
        .c_out(fa_s0_c48_n196_c)
    );

    fa fa_s0_c48_n197 (
        .a(stage0_col48[15]),
        .b(stage0_col48[16]),
        .c_in(stage0_col48[17]),
        .s(fa_s0_c48_n197_s),
        .c_out(fa_s0_c48_n197_c)
    );

    fa fa_s0_c48_n198 (
        .a(stage0_col48[18]),
        .b(stage0_col48[19]),
        .c_in(stage0_col48[20]),
        .s(fa_s0_c48_n198_s),
        .c_out(fa_s0_c48_n198_c)
    );

    fa fa_s0_c48_n199 (
        .a(stage0_col48[21]),
        .b(stage0_col48[22]),
        .c_in(stage0_col48[23]),
        .s(fa_s0_c48_n199_s),
        .c_out(fa_s0_c48_n199_c)
    );

    fa fa_s0_c49_n200 (
        .a(stage0_col49[0]),
        .b(stage0_col49[1]),
        .c_in(stage0_col49[2]),
        .s(fa_s0_c49_n200_s),
        .c_out(fa_s0_c49_n200_c)
    );

    fa fa_s0_c49_n201 (
        .a(stage0_col49[3]),
        .b(stage0_col49[4]),
        .c_in(stage0_col49[5]),
        .s(fa_s0_c49_n201_s),
        .c_out(fa_s0_c49_n201_c)
    );

    fa fa_s0_c49_n202 (
        .a(stage0_col49[6]),
        .b(stage0_col49[7]),
        .c_in(stage0_col49[8]),
        .s(fa_s0_c49_n202_s),
        .c_out(fa_s0_c49_n202_c)
    );

    fa fa_s0_c49_n203 (
        .a(stage0_col49[9]),
        .b(stage0_col49[10]),
        .c_in(stage0_col49[11]),
        .s(fa_s0_c49_n203_s),
        .c_out(fa_s0_c49_n203_c)
    );

    fa fa_s0_c49_n204 (
        .a(stage0_col49[12]),
        .b(stage0_col49[13]),
        .c_in(stage0_col49[14]),
        .s(fa_s0_c49_n204_s),
        .c_out(fa_s0_c49_n204_c)
    );

    fa fa_s0_c49_n205 (
        .a(stage0_col49[15]),
        .b(stage0_col49[16]),
        .c_in(stage0_col49[17]),
        .s(fa_s0_c49_n205_s),
        .c_out(fa_s0_c49_n205_c)
    );

    fa fa_s0_c49_n206 (
        .a(stage0_col49[18]),
        .b(stage0_col49[19]),
        .c_in(stage0_col49[20]),
        .s(fa_s0_c49_n206_s),
        .c_out(fa_s0_c49_n206_c)
    );

    fa fa_s0_c49_n207 (
        .a(stage0_col49[21]),
        .b(stage0_col49[22]),
        .c_in(stage0_col49[23]),
        .s(fa_s0_c49_n207_s),
        .c_out(fa_s0_c49_n207_c)
    );

    fa fa_s0_c50_n208 (
        .a(stage0_col50[0]),
        .b(stage0_col50[1]),
        .c_in(stage0_col50[2]),
        .s(fa_s0_c50_n208_s),
        .c_out(fa_s0_c50_n208_c)
    );

    fa fa_s0_c50_n209 (
        .a(stage0_col50[3]),
        .b(stage0_col50[4]),
        .c_in(stage0_col50[5]),
        .s(fa_s0_c50_n209_s),
        .c_out(fa_s0_c50_n209_c)
    );

    fa fa_s0_c50_n210 (
        .a(stage0_col50[6]),
        .b(stage0_col50[7]),
        .c_in(stage0_col50[8]),
        .s(fa_s0_c50_n210_s),
        .c_out(fa_s0_c50_n210_c)
    );

    fa fa_s0_c50_n211 (
        .a(stage0_col50[9]),
        .b(stage0_col50[10]),
        .c_in(stage0_col50[11]),
        .s(fa_s0_c50_n211_s),
        .c_out(fa_s0_c50_n211_c)
    );

    fa fa_s0_c50_n212 (
        .a(stage0_col50[12]),
        .b(stage0_col50[13]),
        .c_in(stage0_col50[14]),
        .s(fa_s0_c50_n212_s),
        .c_out(fa_s0_c50_n212_c)
    );

    fa fa_s0_c50_n213 (
        .a(stage0_col50[15]),
        .b(stage0_col50[16]),
        .c_in(stage0_col50[17]),
        .s(fa_s0_c50_n213_s),
        .c_out(fa_s0_c50_n213_c)
    );

    fa fa_s0_c50_n214 (
        .a(stage0_col50[18]),
        .b(stage0_col50[19]),
        .c_in(stage0_col50[20]),
        .s(fa_s0_c50_n214_s),
        .c_out(fa_s0_c50_n214_c)
    );

    fa fa_s0_c50_n215 (
        .a(stage0_col50[21]),
        .b(stage0_col50[22]),
        .c_in(stage0_col50[23]),
        .s(fa_s0_c50_n215_s),
        .c_out(fa_s0_c50_n215_c)
    );

    fa fa_s0_c50_n216 (
        .a(stage0_col50[24]),
        .b(stage0_col50[25]),
        .c_in(stage0_col50[26]),
        .s(fa_s0_c50_n216_s),
        .c_out(fa_s0_c50_n216_c)
    );

    fa fa_s0_c51_n217 (
        .a(stage0_col51[0]),
        .b(stage0_col51[1]),
        .c_in(stage0_col51[2]),
        .s(fa_s0_c51_n217_s),
        .c_out(fa_s0_c51_n217_c)
    );

    fa fa_s0_c51_n218 (
        .a(stage0_col51[3]),
        .b(stage0_col51[4]),
        .c_in(stage0_col51[5]),
        .s(fa_s0_c51_n218_s),
        .c_out(fa_s0_c51_n218_c)
    );

    fa fa_s0_c51_n219 (
        .a(stage0_col51[6]),
        .b(stage0_col51[7]),
        .c_in(stage0_col51[8]),
        .s(fa_s0_c51_n219_s),
        .c_out(fa_s0_c51_n219_c)
    );

    fa fa_s0_c51_n220 (
        .a(stage0_col51[9]),
        .b(stage0_col51[10]),
        .c_in(stage0_col51[11]),
        .s(fa_s0_c51_n220_s),
        .c_out(fa_s0_c51_n220_c)
    );

    fa fa_s0_c51_n221 (
        .a(stage0_col51[12]),
        .b(stage0_col51[13]),
        .c_in(stage0_col51[14]),
        .s(fa_s0_c51_n221_s),
        .c_out(fa_s0_c51_n221_c)
    );

    fa fa_s0_c51_n222 (
        .a(stage0_col51[15]),
        .b(stage0_col51[16]),
        .c_in(stage0_col51[17]),
        .s(fa_s0_c51_n222_s),
        .c_out(fa_s0_c51_n222_c)
    );

    fa fa_s0_c51_n223 (
        .a(stage0_col51[18]),
        .b(stage0_col51[19]),
        .c_in(stage0_col51[20]),
        .s(fa_s0_c51_n223_s),
        .c_out(fa_s0_c51_n223_c)
    );

    fa fa_s0_c51_n224 (
        .a(stage0_col51[21]),
        .b(stage0_col51[22]),
        .c_in(stage0_col51[23]),
        .s(fa_s0_c51_n224_s),
        .c_out(fa_s0_c51_n224_c)
    );

    fa fa_s0_c52_n225 (
        .a(stage0_col52[0]),
        .b(stage0_col52[1]),
        .c_in(stage0_col52[2]),
        .s(fa_s0_c52_n225_s),
        .c_out(fa_s0_c52_n225_c)
    );

    fa fa_s0_c52_n226 (
        .a(stage0_col52[3]),
        .b(stage0_col52[4]),
        .c_in(stage0_col52[5]),
        .s(fa_s0_c52_n226_s),
        .c_out(fa_s0_c52_n226_c)
    );

    fa fa_s0_c52_n227 (
        .a(stage0_col52[6]),
        .b(stage0_col52[7]),
        .c_in(stage0_col52[8]),
        .s(fa_s0_c52_n227_s),
        .c_out(fa_s0_c52_n227_c)
    );

    fa fa_s0_c52_n228 (
        .a(stage0_col52[9]),
        .b(stage0_col52[10]),
        .c_in(stage0_col52[11]),
        .s(fa_s0_c52_n228_s),
        .c_out(fa_s0_c52_n228_c)
    );

    fa fa_s0_c52_n229 (
        .a(stage0_col52[12]),
        .b(stage0_col52[13]),
        .c_in(stage0_col52[14]),
        .s(fa_s0_c52_n229_s),
        .c_out(fa_s0_c52_n229_c)
    );

    fa fa_s0_c52_n230 (
        .a(stage0_col52[15]),
        .b(stage0_col52[16]),
        .c_in(stage0_col52[17]),
        .s(fa_s0_c52_n230_s),
        .c_out(fa_s0_c52_n230_c)
    );

    fa fa_s0_c52_n231 (
        .a(stage0_col52[18]),
        .b(stage0_col52[19]),
        .c_in(stage0_col52[20]),
        .s(fa_s0_c52_n231_s),
        .c_out(fa_s0_c52_n231_c)
    );

    fa fa_s0_c52_n232 (
        .a(stage0_col52[21]),
        .b(stage0_col52[22]),
        .c_in(stage0_col52[23]),
        .s(fa_s0_c52_n232_s),
        .c_out(fa_s0_c52_n232_c)
    );

    fa fa_s0_c52_n233 (
        .a(stage0_col52[24]),
        .b(stage0_col52[25]),
        .c_in(stage0_col52[26]),
        .s(fa_s0_c52_n233_s),
        .c_out(fa_s0_c52_n233_c)
    );

    fa fa_s0_c53_n234 (
        .a(stage0_col53[0]),
        .b(stage0_col53[1]),
        .c_in(stage0_col53[2]),
        .s(fa_s0_c53_n234_s),
        .c_out(fa_s0_c53_n234_c)
    );

    fa fa_s0_c53_n235 (
        .a(stage0_col53[3]),
        .b(stage0_col53[4]),
        .c_in(stage0_col53[5]),
        .s(fa_s0_c53_n235_s),
        .c_out(fa_s0_c53_n235_c)
    );

    fa fa_s0_c53_n236 (
        .a(stage0_col53[6]),
        .b(stage0_col53[7]),
        .c_in(stage0_col53[8]),
        .s(fa_s0_c53_n236_s),
        .c_out(fa_s0_c53_n236_c)
    );

    fa fa_s0_c53_n237 (
        .a(stage0_col53[9]),
        .b(stage0_col53[10]),
        .c_in(stage0_col53[11]),
        .s(fa_s0_c53_n237_s),
        .c_out(fa_s0_c53_n237_c)
    );

    fa fa_s0_c53_n238 (
        .a(stage0_col53[12]),
        .b(stage0_col53[13]),
        .c_in(stage0_col53[14]),
        .s(fa_s0_c53_n238_s),
        .c_out(fa_s0_c53_n238_c)
    );

    fa fa_s0_c53_n239 (
        .a(stage0_col53[15]),
        .b(stage0_col53[16]),
        .c_in(stage0_col53[17]),
        .s(fa_s0_c53_n239_s),
        .c_out(fa_s0_c53_n239_c)
    );

    fa fa_s0_c53_n240 (
        .a(stage0_col53[18]),
        .b(stage0_col53[19]),
        .c_in(stage0_col53[20]),
        .s(fa_s0_c53_n240_s),
        .c_out(fa_s0_c53_n240_c)
    );

    fa fa_s0_c53_n241 (
        .a(stage0_col53[21]),
        .b(stage0_col53[22]),
        .c_in(stage0_col53[23]),
        .s(fa_s0_c53_n241_s),
        .c_out(fa_s0_c53_n241_c)
    );

    fa fa_s0_c53_n242 (
        .a(stage0_col53[24]),
        .b(stage0_col53[25]),
        .c_in(stage0_col53[26]),
        .s(fa_s0_c53_n242_s),
        .c_out(fa_s0_c53_n242_c)
    );

    fa fa_s0_c54_n243 (
        .a(stage0_col54[0]),
        .b(stage0_col54[1]),
        .c_in(stage0_col54[2]),
        .s(fa_s0_c54_n243_s),
        .c_out(fa_s0_c54_n243_c)
    );

    fa fa_s0_c54_n244 (
        .a(stage0_col54[3]),
        .b(stage0_col54[4]),
        .c_in(stage0_col54[5]),
        .s(fa_s0_c54_n244_s),
        .c_out(fa_s0_c54_n244_c)
    );

    fa fa_s0_c54_n245 (
        .a(stage0_col54[6]),
        .b(stage0_col54[7]),
        .c_in(stage0_col54[8]),
        .s(fa_s0_c54_n245_s),
        .c_out(fa_s0_c54_n245_c)
    );

    fa fa_s0_c54_n246 (
        .a(stage0_col54[9]),
        .b(stage0_col54[10]),
        .c_in(stage0_col54[11]),
        .s(fa_s0_c54_n246_s),
        .c_out(fa_s0_c54_n246_c)
    );

    fa fa_s0_c54_n247 (
        .a(stage0_col54[12]),
        .b(stage0_col54[13]),
        .c_in(stage0_col54[14]),
        .s(fa_s0_c54_n247_s),
        .c_out(fa_s0_c54_n247_c)
    );

    fa fa_s0_c54_n248 (
        .a(stage0_col54[15]),
        .b(stage0_col54[16]),
        .c_in(stage0_col54[17]),
        .s(fa_s0_c54_n248_s),
        .c_out(fa_s0_c54_n248_c)
    );

    fa fa_s0_c54_n249 (
        .a(stage0_col54[18]),
        .b(stage0_col54[19]),
        .c_in(stage0_col54[20]),
        .s(fa_s0_c54_n249_s),
        .c_out(fa_s0_c54_n249_c)
    );

    fa fa_s0_c54_n250 (
        .a(stage0_col54[21]),
        .b(stage0_col54[22]),
        .c_in(stage0_col54[23]),
        .s(fa_s0_c54_n250_s),
        .c_out(fa_s0_c54_n250_c)
    );

    fa fa_s0_c54_n251 (
        .a(stage0_col54[24]),
        .b(stage0_col54[25]),
        .c_in(stage0_col54[26]),
        .s(fa_s0_c54_n251_s),
        .c_out(fa_s0_c54_n251_c)
    );

    fa fa_s0_c55_n252 (
        .a(stage0_col55[0]),
        .b(stage0_col55[1]),
        .c_in(stage0_col55[2]),
        .s(fa_s0_c55_n252_s),
        .c_out(fa_s0_c55_n252_c)
    );

    fa fa_s0_c55_n253 (
        .a(stage0_col55[3]),
        .b(stage0_col55[4]),
        .c_in(stage0_col55[5]),
        .s(fa_s0_c55_n253_s),
        .c_out(fa_s0_c55_n253_c)
    );

    fa fa_s0_c55_n254 (
        .a(stage0_col55[6]),
        .b(stage0_col55[7]),
        .c_in(stage0_col55[8]),
        .s(fa_s0_c55_n254_s),
        .c_out(fa_s0_c55_n254_c)
    );

    fa fa_s0_c55_n255 (
        .a(stage0_col55[9]),
        .b(stage0_col55[10]),
        .c_in(stage0_col55[11]),
        .s(fa_s0_c55_n255_s),
        .c_out(fa_s0_c55_n255_c)
    );

    fa fa_s0_c55_n256 (
        .a(stage0_col55[12]),
        .b(stage0_col55[13]),
        .c_in(stage0_col55[14]),
        .s(fa_s0_c55_n256_s),
        .c_out(fa_s0_c55_n256_c)
    );

    fa fa_s0_c55_n257 (
        .a(stage0_col55[15]),
        .b(stage0_col55[16]),
        .c_in(stage0_col55[17]),
        .s(fa_s0_c55_n257_s),
        .c_out(fa_s0_c55_n257_c)
    );

    fa fa_s0_c55_n258 (
        .a(stage0_col55[18]),
        .b(stage0_col55[19]),
        .c_in(stage0_col55[20]),
        .s(fa_s0_c55_n258_s),
        .c_out(fa_s0_c55_n258_c)
    );

    fa fa_s0_c55_n259 (
        .a(stage0_col55[21]),
        .b(stage0_col55[22]),
        .c_in(stage0_col55[23]),
        .s(fa_s0_c55_n259_s),
        .c_out(fa_s0_c55_n259_c)
    );

    fa fa_s0_c55_n260 (
        .a(stage0_col55[24]),
        .b(stage0_col55[25]),
        .c_in(stage0_col55[26]),
        .s(fa_s0_c55_n260_s),
        .c_out(fa_s0_c55_n260_c)
    );

    fa fa_s0_c56_n261 (
        .a(stage0_col56[0]),
        .b(stage0_col56[1]),
        .c_in(stage0_col56[2]),
        .s(fa_s0_c56_n261_s),
        .c_out(fa_s0_c56_n261_c)
    );

    fa fa_s0_c56_n262 (
        .a(stage0_col56[3]),
        .b(stage0_col56[4]),
        .c_in(stage0_col56[5]),
        .s(fa_s0_c56_n262_s),
        .c_out(fa_s0_c56_n262_c)
    );

    fa fa_s0_c56_n263 (
        .a(stage0_col56[6]),
        .b(stage0_col56[7]),
        .c_in(stage0_col56[8]),
        .s(fa_s0_c56_n263_s),
        .c_out(fa_s0_c56_n263_c)
    );

    fa fa_s0_c56_n264 (
        .a(stage0_col56[9]),
        .b(stage0_col56[10]),
        .c_in(stage0_col56[11]),
        .s(fa_s0_c56_n264_s),
        .c_out(fa_s0_c56_n264_c)
    );

    fa fa_s0_c56_n265 (
        .a(stage0_col56[12]),
        .b(stage0_col56[13]),
        .c_in(stage0_col56[14]),
        .s(fa_s0_c56_n265_s),
        .c_out(fa_s0_c56_n265_c)
    );

    fa fa_s0_c56_n266 (
        .a(stage0_col56[15]),
        .b(stage0_col56[16]),
        .c_in(stage0_col56[17]),
        .s(fa_s0_c56_n266_s),
        .c_out(fa_s0_c56_n266_c)
    );

    fa fa_s0_c56_n267 (
        .a(stage0_col56[18]),
        .b(stage0_col56[19]),
        .c_in(stage0_col56[20]),
        .s(fa_s0_c56_n267_s),
        .c_out(fa_s0_c56_n267_c)
    );

    fa fa_s0_c56_n268 (
        .a(stage0_col56[21]),
        .b(stage0_col56[22]),
        .c_in(stage0_col56[23]),
        .s(fa_s0_c56_n268_s),
        .c_out(fa_s0_c56_n268_c)
    );

    fa fa_s0_c56_n269 (
        .a(stage0_col56[24]),
        .b(stage0_col56[25]),
        .c_in(stage0_col56[26]),
        .s(fa_s0_c56_n269_s),
        .c_out(fa_s0_c56_n269_c)
    );

    fa fa_s0_c56_n270 (
        .a(stage0_col56[27]),
        .b(stage0_col56[28]),
        .c_in(stage0_col56[29]),
        .s(fa_s0_c56_n270_s),
        .c_out(fa_s0_c56_n270_c)
    );

    fa fa_s0_c57_n271 (
        .a(stage0_col57[0]),
        .b(stage0_col57[1]),
        .c_in(stage0_col57[2]),
        .s(fa_s0_c57_n271_s),
        .c_out(fa_s0_c57_n271_c)
    );

    fa fa_s0_c57_n272 (
        .a(stage0_col57[3]),
        .b(stage0_col57[4]),
        .c_in(stage0_col57[5]),
        .s(fa_s0_c57_n272_s),
        .c_out(fa_s0_c57_n272_c)
    );

    fa fa_s0_c57_n273 (
        .a(stage0_col57[6]),
        .b(stage0_col57[7]),
        .c_in(stage0_col57[8]),
        .s(fa_s0_c57_n273_s),
        .c_out(fa_s0_c57_n273_c)
    );

    fa fa_s0_c57_n274 (
        .a(stage0_col57[9]),
        .b(stage0_col57[10]),
        .c_in(stage0_col57[11]),
        .s(fa_s0_c57_n274_s),
        .c_out(fa_s0_c57_n274_c)
    );

    fa fa_s0_c57_n275 (
        .a(stage0_col57[12]),
        .b(stage0_col57[13]),
        .c_in(stage0_col57[14]),
        .s(fa_s0_c57_n275_s),
        .c_out(fa_s0_c57_n275_c)
    );

    fa fa_s0_c57_n276 (
        .a(stage0_col57[15]),
        .b(stage0_col57[16]),
        .c_in(stage0_col57[17]),
        .s(fa_s0_c57_n276_s),
        .c_out(fa_s0_c57_n276_c)
    );

    fa fa_s0_c57_n277 (
        .a(stage0_col57[18]),
        .b(stage0_col57[19]),
        .c_in(stage0_col57[20]),
        .s(fa_s0_c57_n277_s),
        .c_out(fa_s0_c57_n277_c)
    );

    fa fa_s0_c57_n278 (
        .a(stage0_col57[21]),
        .b(stage0_col57[22]),
        .c_in(stage0_col57[23]),
        .s(fa_s0_c57_n278_s),
        .c_out(fa_s0_c57_n278_c)
    );

    fa fa_s0_c57_n279 (
        .a(stage0_col57[24]),
        .b(stage0_col57[25]),
        .c_in(stage0_col57[26]),
        .s(fa_s0_c57_n279_s),
        .c_out(fa_s0_c57_n279_c)
    );

    fa fa_s0_c58_n280 (
        .a(stage0_col58[0]),
        .b(stage0_col58[1]),
        .c_in(stage0_col58[2]),
        .s(fa_s0_c58_n280_s),
        .c_out(fa_s0_c58_n280_c)
    );

    fa fa_s0_c58_n281 (
        .a(stage0_col58[3]),
        .b(stage0_col58[4]),
        .c_in(stage0_col58[5]),
        .s(fa_s0_c58_n281_s),
        .c_out(fa_s0_c58_n281_c)
    );

    fa fa_s0_c58_n282 (
        .a(stage0_col58[6]),
        .b(stage0_col58[7]),
        .c_in(stage0_col58[8]),
        .s(fa_s0_c58_n282_s),
        .c_out(fa_s0_c58_n282_c)
    );

    fa fa_s0_c58_n283 (
        .a(stage0_col58[9]),
        .b(stage0_col58[10]),
        .c_in(stage0_col58[11]),
        .s(fa_s0_c58_n283_s),
        .c_out(fa_s0_c58_n283_c)
    );

    fa fa_s0_c58_n284 (
        .a(stage0_col58[12]),
        .b(stage0_col58[13]),
        .c_in(stage0_col58[14]),
        .s(fa_s0_c58_n284_s),
        .c_out(fa_s0_c58_n284_c)
    );

    fa fa_s0_c58_n285 (
        .a(stage0_col58[15]),
        .b(stage0_col58[16]),
        .c_in(stage0_col58[17]),
        .s(fa_s0_c58_n285_s),
        .c_out(fa_s0_c58_n285_c)
    );

    fa fa_s0_c58_n286 (
        .a(stage0_col58[18]),
        .b(stage0_col58[19]),
        .c_in(stage0_col58[20]),
        .s(fa_s0_c58_n286_s),
        .c_out(fa_s0_c58_n286_c)
    );

    fa fa_s0_c58_n287 (
        .a(stage0_col58[21]),
        .b(stage0_col58[22]),
        .c_in(stage0_col58[23]),
        .s(fa_s0_c58_n287_s),
        .c_out(fa_s0_c58_n287_c)
    );

    fa fa_s0_c58_n288 (
        .a(stage0_col58[24]),
        .b(stage0_col58[25]),
        .c_in(stage0_col58[26]),
        .s(fa_s0_c58_n288_s),
        .c_out(fa_s0_c58_n288_c)
    );

    fa fa_s0_c58_n289 (
        .a(stage0_col58[27]),
        .b(stage0_col58[28]),
        .c_in(stage0_col58[29]),
        .s(fa_s0_c58_n289_s),
        .c_out(fa_s0_c58_n289_c)
    );

    fa fa_s0_c59_n290 (
        .a(stage0_col59[0]),
        .b(stage0_col59[1]),
        .c_in(stage0_col59[2]),
        .s(fa_s0_c59_n290_s),
        .c_out(fa_s0_c59_n290_c)
    );

    fa fa_s0_c59_n291 (
        .a(stage0_col59[3]),
        .b(stage0_col59[4]),
        .c_in(stage0_col59[5]),
        .s(fa_s0_c59_n291_s),
        .c_out(fa_s0_c59_n291_c)
    );

    fa fa_s0_c59_n292 (
        .a(stage0_col59[6]),
        .b(stage0_col59[7]),
        .c_in(stage0_col59[8]),
        .s(fa_s0_c59_n292_s),
        .c_out(fa_s0_c59_n292_c)
    );

    fa fa_s0_c59_n293 (
        .a(stage0_col59[9]),
        .b(stage0_col59[10]),
        .c_in(stage0_col59[11]),
        .s(fa_s0_c59_n293_s),
        .c_out(fa_s0_c59_n293_c)
    );

    fa fa_s0_c59_n294 (
        .a(stage0_col59[12]),
        .b(stage0_col59[13]),
        .c_in(stage0_col59[14]),
        .s(fa_s0_c59_n294_s),
        .c_out(fa_s0_c59_n294_c)
    );

    fa fa_s0_c59_n295 (
        .a(stage0_col59[15]),
        .b(stage0_col59[16]),
        .c_in(stage0_col59[17]),
        .s(fa_s0_c59_n295_s),
        .c_out(fa_s0_c59_n295_c)
    );

    fa fa_s0_c59_n296 (
        .a(stage0_col59[18]),
        .b(stage0_col59[19]),
        .c_in(stage0_col59[20]),
        .s(fa_s0_c59_n296_s),
        .c_out(fa_s0_c59_n296_c)
    );

    fa fa_s0_c59_n297 (
        .a(stage0_col59[21]),
        .b(stage0_col59[22]),
        .c_in(stage0_col59[23]),
        .s(fa_s0_c59_n297_s),
        .c_out(fa_s0_c59_n297_c)
    );

    fa fa_s0_c59_n298 (
        .a(stage0_col59[24]),
        .b(stage0_col59[25]),
        .c_in(stage0_col59[26]),
        .s(fa_s0_c59_n298_s),
        .c_out(fa_s0_c59_n298_c)
    );

    fa fa_s0_c59_n299 (
        .a(stage0_col59[27]),
        .b(stage0_col59[28]),
        .c_in(stage0_col59[29]),
        .s(fa_s0_c59_n299_s),
        .c_out(fa_s0_c59_n299_c)
    );

    fa fa_s0_c60_n300 (
        .a(stage0_col60[0]),
        .b(stage0_col60[1]),
        .c_in(stage0_col60[2]),
        .s(fa_s0_c60_n300_s),
        .c_out(fa_s0_c60_n300_c)
    );

    fa fa_s0_c60_n301 (
        .a(stage0_col60[3]),
        .b(stage0_col60[4]),
        .c_in(stage0_col60[5]),
        .s(fa_s0_c60_n301_s),
        .c_out(fa_s0_c60_n301_c)
    );

    fa fa_s0_c60_n302 (
        .a(stage0_col60[6]),
        .b(stage0_col60[7]),
        .c_in(stage0_col60[8]),
        .s(fa_s0_c60_n302_s),
        .c_out(fa_s0_c60_n302_c)
    );

    fa fa_s0_c60_n303 (
        .a(stage0_col60[9]),
        .b(stage0_col60[10]),
        .c_in(stage0_col60[11]),
        .s(fa_s0_c60_n303_s),
        .c_out(fa_s0_c60_n303_c)
    );

    fa fa_s0_c60_n304 (
        .a(stage0_col60[12]),
        .b(stage0_col60[13]),
        .c_in(stage0_col60[14]),
        .s(fa_s0_c60_n304_s),
        .c_out(fa_s0_c60_n304_c)
    );

    fa fa_s0_c60_n305 (
        .a(stage0_col60[15]),
        .b(stage0_col60[16]),
        .c_in(stage0_col60[17]),
        .s(fa_s0_c60_n305_s),
        .c_out(fa_s0_c60_n305_c)
    );

    fa fa_s0_c60_n306 (
        .a(stage0_col60[18]),
        .b(stage0_col60[19]),
        .c_in(stage0_col60[20]),
        .s(fa_s0_c60_n306_s),
        .c_out(fa_s0_c60_n306_c)
    );

    fa fa_s0_c60_n307 (
        .a(stage0_col60[21]),
        .b(stage0_col60[22]),
        .c_in(stage0_col60[23]),
        .s(fa_s0_c60_n307_s),
        .c_out(fa_s0_c60_n307_c)
    );

    fa fa_s0_c60_n308 (
        .a(stage0_col60[24]),
        .b(stage0_col60[25]),
        .c_in(stage0_col60[26]),
        .s(fa_s0_c60_n308_s),
        .c_out(fa_s0_c60_n308_c)
    );

    fa fa_s0_c60_n309 (
        .a(stage0_col60[27]),
        .b(stage0_col60[28]),
        .c_in(stage0_col60[29]),
        .s(fa_s0_c60_n309_s),
        .c_out(fa_s0_c60_n309_c)
    );

    fa fa_s0_c61_n310 (
        .a(stage0_col61[0]),
        .b(stage0_col61[1]),
        .c_in(stage0_col61[2]),
        .s(fa_s0_c61_n310_s),
        .c_out(fa_s0_c61_n310_c)
    );

    fa fa_s0_c61_n311 (
        .a(stage0_col61[3]),
        .b(stage0_col61[4]),
        .c_in(stage0_col61[5]),
        .s(fa_s0_c61_n311_s),
        .c_out(fa_s0_c61_n311_c)
    );

    fa fa_s0_c61_n312 (
        .a(stage0_col61[6]),
        .b(stage0_col61[7]),
        .c_in(stage0_col61[8]),
        .s(fa_s0_c61_n312_s),
        .c_out(fa_s0_c61_n312_c)
    );

    fa fa_s0_c61_n313 (
        .a(stage0_col61[9]),
        .b(stage0_col61[10]),
        .c_in(stage0_col61[11]),
        .s(fa_s0_c61_n313_s),
        .c_out(fa_s0_c61_n313_c)
    );

    fa fa_s0_c61_n314 (
        .a(stage0_col61[12]),
        .b(stage0_col61[13]),
        .c_in(stage0_col61[14]),
        .s(fa_s0_c61_n314_s),
        .c_out(fa_s0_c61_n314_c)
    );

    fa fa_s0_c61_n315 (
        .a(stage0_col61[15]),
        .b(stage0_col61[16]),
        .c_in(stage0_col61[17]),
        .s(fa_s0_c61_n315_s),
        .c_out(fa_s0_c61_n315_c)
    );

    fa fa_s0_c61_n316 (
        .a(stage0_col61[18]),
        .b(stage0_col61[19]),
        .c_in(stage0_col61[20]),
        .s(fa_s0_c61_n316_s),
        .c_out(fa_s0_c61_n316_c)
    );

    fa fa_s0_c61_n317 (
        .a(stage0_col61[21]),
        .b(stage0_col61[22]),
        .c_in(stage0_col61[23]),
        .s(fa_s0_c61_n317_s),
        .c_out(fa_s0_c61_n317_c)
    );

    fa fa_s0_c61_n318 (
        .a(stage0_col61[24]),
        .b(stage0_col61[25]),
        .c_in(stage0_col61[26]),
        .s(fa_s0_c61_n318_s),
        .c_out(fa_s0_c61_n318_c)
    );

    fa fa_s0_c61_n319 (
        .a(stage0_col61[27]),
        .b(stage0_col61[28]),
        .c_in(stage0_col61[29]),
        .s(fa_s0_c61_n319_s),
        .c_out(fa_s0_c61_n319_c)
    );

    fa fa_s0_c62_n320 (
        .a(stage0_col62[0]),
        .b(stage0_col62[1]),
        .c_in(stage0_col62[2]),
        .s(fa_s0_c62_n320_s),
        .c_out(fa_s0_c62_n320_c)
    );

    fa fa_s0_c62_n321 (
        .a(stage0_col62[3]),
        .b(stage0_col62[4]),
        .c_in(stage0_col62[5]),
        .s(fa_s0_c62_n321_s),
        .c_out(fa_s0_c62_n321_c)
    );

    fa fa_s0_c62_n322 (
        .a(stage0_col62[6]),
        .b(stage0_col62[7]),
        .c_in(stage0_col62[8]),
        .s(fa_s0_c62_n322_s),
        .c_out(fa_s0_c62_n322_c)
    );

    fa fa_s0_c62_n323 (
        .a(stage0_col62[9]),
        .b(stage0_col62[10]),
        .c_in(stage0_col62[11]),
        .s(fa_s0_c62_n323_s),
        .c_out(fa_s0_c62_n323_c)
    );

    fa fa_s0_c62_n324 (
        .a(stage0_col62[12]),
        .b(stage0_col62[13]),
        .c_in(stage0_col62[14]),
        .s(fa_s0_c62_n324_s),
        .c_out(fa_s0_c62_n324_c)
    );

    fa fa_s0_c62_n325 (
        .a(stage0_col62[15]),
        .b(stage0_col62[16]),
        .c_in(stage0_col62[17]),
        .s(fa_s0_c62_n325_s),
        .c_out(fa_s0_c62_n325_c)
    );

    fa fa_s0_c62_n326 (
        .a(stage0_col62[18]),
        .b(stage0_col62[19]),
        .c_in(stage0_col62[20]),
        .s(fa_s0_c62_n326_s),
        .c_out(fa_s0_c62_n326_c)
    );

    fa fa_s0_c62_n327 (
        .a(stage0_col62[21]),
        .b(stage0_col62[22]),
        .c_in(stage0_col62[23]),
        .s(fa_s0_c62_n327_s),
        .c_out(fa_s0_c62_n327_c)
    );

    fa fa_s0_c62_n328 (
        .a(stage0_col62[24]),
        .b(stage0_col62[25]),
        .c_in(stage0_col62[26]),
        .s(fa_s0_c62_n328_s),
        .c_out(fa_s0_c62_n328_c)
    );

    fa fa_s0_c62_n329 (
        .a(stage0_col62[27]),
        .b(stage0_col62[28]),
        .c_in(stage0_col62[29]),
        .s(fa_s0_c62_n329_s),
        .c_out(fa_s0_c62_n329_c)
    );

    fa fa_s0_c62_n330 (
        .a(stage0_col62[30]),
        .b(stage0_col62[31]),
        .c_in(stage0_col62[32]),
        .s(fa_s0_c62_n330_s),
        .c_out(fa_s0_c62_n330_c)
    );

    fa fa_s0_c63_n331 (
        .a(stage0_col63[0]),
        .b(stage0_col63[1]),
        .c_in(stage0_col63[2]),
        .s(fa_s0_c63_n331_s),
        .c_out(fa_s0_c63_n331_c)
    );

    fa fa_s0_c63_n332 (
        .a(stage0_col63[3]),
        .b(stage0_col63[4]),
        .c_in(stage0_col63[5]),
        .s(fa_s0_c63_n332_s),
        .c_out(fa_s0_c63_n332_c)
    );

    fa fa_s0_c63_n333 (
        .a(stage0_col63[6]),
        .b(stage0_col63[7]),
        .c_in(stage0_col63[8]),
        .s(fa_s0_c63_n333_s),
        .c_out(fa_s0_c63_n333_c)
    );

    fa fa_s0_c63_n334 (
        .a(stage0_col63[9]),
        .b(stage0_col63[10]),
        .c_in(stage0_col63[11]),
        .s(fa_s0_c63_n334_s),
        .c_out(fa_s0_c63_n334_c)
    );

    fa fa_s0_c63_n335 (
        .a(stage0_col63[12]),
        .b(stage0_col63[13]),
        .c_in(stage0_col63[14]),
        .s(fa_s0_c63_n335_s),
        .c_out(fa_s0_c63_n335_c)
    );

    fa fa_s0_c63_n336 (
        .a(stage0_col63[15]),
        .b(stage0_col63[16]),
        .c_in(stage0_col63[17]),
        .s(fa_s0_c63_n336_s),
        .c_out(fa_s0_c63_n336_c)
    );

    fa fa_s0_c63_n337 (
        .a(stage0_col63[18]),
        .b(stage0_col63[19]),
        .c_in(stage0_col63[20]),
        .s(fa_s0_c63_n337_s),
        .c_out(fa_s0_c63_n337_c)
    );

    fa fa_s0_c63_n338 (
        .a(stage0_col63[21]),
        .b(stage0_col63[22]),
        .c_in(stage0_col63[23]),
        .s(fa_s0_c63_n338_s),
        .c_out(fa_s0_c63_n338_c)
    );

    fa fa_s0_c63_n339 (
        .a(stage0_col63[24]),
        .b(stage0_col63[25]),
        .c_in(stage0_col63[26]),
        .s(fa_s0_c63_n339_s),
        .c_out(fa_s0_c63_n339_c)
    );

    fa fa_s0_c63_n340 (
        .a(stage0_col63[27]),
        .b(stage0_col63[28]),
        .c_in(stage0_col63[29]),
        .s(fa_s0_c63_n340_s),
        .c_out(fa_s0_c63_n340_c)
    );

    fa fa_s0_c64_n341 (
        .a(stage0_col64[0]),
        .b(stage0_col64[1]),
        .c_in(stage0_col64[2]),
        .s(fa_s0_c64_n341_s),
        .c_out(fa_s0_c64_n341_c)
    );

    fa fa_s0_c64_n342 (
        .a(stage0_col64[3]),
        .b(stage0_col64[4]),
        .c_in(stage0_col64[5]),
        .s(fa_s0_c64_n342_s),
        .c_out(fa_s0_c64_n342_c)
    );

    fa fa_s0_c64_n343 (
        .a(stage0_col64[6]),
        .b(stage0_col64[7]),
        .c_in(stage0_col64[8]),
        .s(fa_s0_c64_n343_s),
        .c_out(fa_s0_c64_n343_c)
    );

    fa fa_s0_c64_n344 (
        .a(stage0_col64[9]),
        .b(stage0_col64[10]),
        .c_in(stage0_col64[11]),
        .s(fa_s0_c64_n344_s),
        .c_out(fa_s0_c64_n344_c)
    );

    fa fa_s0_c64_n345 (
        .a(stage0_col64[12]),
        .b(stage0_col64[13]),
        .c_in(stage0_col64[14]),
        .s(fa_s0_c64_n345_s),
        .c_out(fa_s0_c64_n345_c)
    );

    fa fa_s0_c64_n346 (
        .a(stage0_col64[15]),
        .b(stage0_col64[16]),
        .c_in(stage0_col64[17]),
        .s(fa_s0_c64_n346_s),
        .c_out(fa_s0_c64_n346_c)
    );

    fa fa_s0_c64_n347 (
        .a(stage0_col64[18]),
        .b(stage0_col64[19]),
        .c_in(stage0_col64[20]),
        .s(fa_s0_c64_n347_s),
        .c_out(fa_s0_c64_n347_c)
    );

    fa fa_s0_c64_n348 (
        .a(stage0_col64[21]),
        .b(stage0_col64[22]),
        .c_in(stage0_col64[23]),
        .s(fa_s0_c64_n348_s),
        .c_out(fa_s0_c64_n348_c)
    );

    fa fa_s0_c64_n349 (
        .a(stage0_col64[24]),
        .b(stage0_col64[25]),
        .c_in(stage0_col64[26]),
        .s(fa_s0_c64_n349_s),
        .c_out(fa_s0_c64_n349_c)
    );

    fa fa_s0_c64_n350 (
        .a(stage0_col64[27]),
        .b(stage0_col64[28]),
        .c_in(stage0_col64[29]),
        .s(fa_s0_c64_n350_s),
        .c_out(fa_s0_c64_n350_c)
    );

    fa fa_s0_c64_n351 (
        .a(stage0_col64[30]),
        .b(stage0_col64[31]),
        .c_in(stage0_col64[32]),
        .s(fa_s0_c64_n351_s),
        .c_out(fa_s0_c64_n351_c)
    );

    fa fa_s0_c65_n352 (
        .a(stage0_col65[0]),
        .b(stage0_col65[1]),
        .c_in(stage0_col65[2]),
        .s(fa_s0_c65_n352_s),
        .c_out(fa_s0_c65_n352_c)
    );

    fa fa_s0_c65_n353 (
        .a(stage0_col65[3]),
        .b(stage0_col65[4]),
        .c_in(stage0_col65[5]),
        .s(fa_s0_c65_n353_s),
        .c_out(fa_s0_c65_n353_c)
    );

    fa fa_s0_c65_n354 (
        .a(stage0_col65[6]),
        .b(stage0_col65[7]),
        .c_in(stage0_col65[8]),
        .s(fa_s0_c65_n354_s),
        .c_out(fa_s0_c65_n354_c)
    );

    fa fa_s0_c65_n355 (
        .a(stage0_col65[9]),
        .b(stage0_col65[10]),
        .c_in(stage0_col65[11]),
        .s(fa_s0_c65_n355_s),
        .c_out(fa_s0_c65_n355_c)
    );

    fa fa_s0_c65_n356 (
        .a(stage0_col65[12]),
        .b(stage0_col65[13]),
        .c_in(stage0_col65[14]),
        .s(fa_s0_c65_n356_s),
        .c_out(fa_s0_c65_n356_c)
    );

    fa fa_s0_c65_n357 (
        .a(stage0_col65[15]),
        .b(stage0_col65[16]),
        .c_in(stage0_col65[17]),
        .s(fa_s0_c65_n357_s),
        .c_out(fa_s0_c65_n357_c)
    );

    fa fa_s0_c65_n358 (
        .a(stage0_col65[18]),
        .b(stage0_col65[19]),
        .c_in(stage0_col65[20]),
        .s(fa_s0_c65_n358_s),
        .c_out(fa_s0_c65_n358_c)
    );

    fa fa_s0_c65_n359 (
        .a(stage0_col65[21]),
        .b(stage0_col65[22]),
        .c_in(stage0_col65[23]),
        .s(fa_s0_c65_n359_s),
        .c_out(fa_s0_c65_n359_c)
    );

    fa fa_s0_c65_n360 (
        .a(stage0_col65[24]),
        .b(stage0_col65[25]),
        .c_in(stage0_col65[26]),
        .s(fa_s0_c65_n360_s),
        .c_out(fa_s0_c65_n360_c)
    );

    fa fa_s0_c65_n361 (
        .a(stage0_col65[27]),
        .b(stage0_col65[28]),
        .c_in(stage0_col65[29]),
        .s(fa_s0_c65_n361_s),
        .c_out(fa_s0_c65_n361_c)
    );

    fa fa_s0_c66_n362 (
        .a(stage0_col66[0]),
        .b(stage0_col66[1]),
        .c_in(stage0_col66[2]),
        .s(fa_s0_c66_n362_s),
        .c_out(fa_s0_c66_n362_c)
    );

    fa fa_s0_c66_n363 (
        .a(stage0_col66[3]),
        .b(stage0_col66[4]),
        .c_in(stage0_col66[5]),
        .s(fa_s0_c66_n363_s),
        .c_out(fa_s0_c66_n363_c)
    );

    fa fa_s0_c66_n364 (
        .a(stage0_col66[6]),
        .b(stage0_col66[7]),
        .c_in(stage0_col66[8]),
        .s(fa_s0_c66_n364_s),
        .c_out(fa_s0_c66_n364_c)
    );

    fa fa_s0_c66_n365 (
        .a(stage0_col66[9]),
        .b(stage0_col66[10]),
        .c_in(stage0_col66[11]),
        .s(fa_s0_c66_n365_s),
        .c_out(fa_s0_c66_n365_c)
    );

    fa fa_s0_c66_n366 (
        .a(stage0_col66[12]),
        .b(stage0_col66[13]),
        .c_in(stage0_col66[14]),
        .s(fa_s0_c66_n366_s),
        .c_out(fa_s0_c66_n366_c)
    );

    fa fa_s0_c66_n367 (
        .a(stage0_col66[15]),
        .b(stage0_col66[16]),
        .c_in(stage0_col66[17]),
        .s(fa_s0_c66_n367_s),
        .c_out(fa_s0_c66_n367_c)
    );

    fa fa_s0_c66_n368 (
        .a(stage0_col66[18]),
        .b(stage0_col66[19]),
        .c_in(stage0_col66[20]),
        .s(fa_s0_c66_n368_s),
        .c_out(fa_s0_c66_n368_c)
    );

    fa fa_s0_c66_n369 (
        .a(stage0_col66[21]),
        .b(stage0_col66[22]),
        .c_in(stage0_col66[23]),
        .s(fa_s0_c66_n369_s),
        .c_out(fa_s0_c66_n369_c)
    );

    fa fa_s0_c66_n370 (
        .a(stage0_col66[24]),
        .b(stage0_col66[25]),
        .c_in(stage0_col66[26]),
        .s(fa_s0_c66_n370_s),
        .c_out(fa_s0_c66_n370_c)
    );

    fa fa_s0_c66_n371 (
        .a(stage0_col66[27]),
        .b(stage0_col66[28]),
        .c_in(stage0_col66[29]),
        .s(fa_s0_c66_n371_s),
        .c_out(fa_s0_c66_n371_c)
    );

    fa fa_s0_c66_n372 (
        .a(stage0_col66[30]),
        .b(stage0_col66[31]),
        .c_in(stage0_col66[32]),
        .s(fa_s0_c66_n372_s),
        .c_out(fa_s0_c66_n372_c)
    );

    fa fa_s0_c67_n373 (
        .a(stage0_col67[0]),
        .b(stage0_col67[1]),
        .c_in(stage0_col67[2]),
        .s(fa_s0_c67_n373_s),
        .c_out(fa_s0_c67_n373_c)
    );

    fa fa_s0_c67_n374 (
        .a(stage0_col67[3]),
        .b(stage0_col67[4]),
        .c_in(stage0_col67[5]),
        .s(fa_s0_c67_n374_s),
        .c_out(fa_s0_c67_n374_c)
    );

    fa fa_s0_c67_n375 (
        .a(stage0_col67[6]),
        .b(stage0_col67[7]),
        .c_in(stage0_col67[8]),
        .s(fa_s0_c67_n375_s),
        .c_out(fa_s0_c67_n375_c)
    );

    fa fa_s0_c67_n376 (
        .a(stage0_col67[9]),
        .b(stage0_col67[10]),
        .c_in(stage0_col67[11]),
        .s(fa_s0_c67_n376_s),
        .c_out(fa_s0_c67_n376_c)
    );

    fa fa_s0_c67_n377 (
        .a(stage0_col67[12]),
        .b(stage0_col67[13]),
        .c_in(stage0_col67[14]),
        .s(fa_s0_c67_n377_s),
        .c_out(fa_s0_c67_n377_c)
    );

    fa fa_s0_c67_n378 (
        .a(stage0_col67[15]),
        .b(stage0_col67[16]),
        .c_in(stage0_col67[17]),
        .s(fa_s0_c67_n378_s),
        .c_out(fa_s0_c67_n378_c)
    );

    fa fa_s0_c67_n379 (
        .a(stage0_col67[18]),
        .b(stage0_col67[19]),
        .c_in(stage0_col67[20]),
        .s(fa_s0_c67_n379_s),
        .c_out(fa_s0_c67_n379_c)
    );

    fa fa_s0_c67_n380 (
        .a(stage0_col67[21]),
        .b(stage0_col67[22]),
        .c_in(stage0_col67[23]),
        .s(fa_s0_c67_n380_s),
        .c_out(fa_s0_c67_n380_c)
    );

    fa fa_s0_c67_n381 (
        .a(stage0_col67[24]),
        .b(stage0_col67[25]),
        .c_in(stage0_col67[26]),
        .s(fa_s0_c67_n381_s),
        .c_out(fa_s0_c67_n381_c)
    );

    fa fa_s0_c67_n382 (
        .a(stage0_col67[27]),
        .b(stage0_col67[28]),
        .c_in(stage0_col67[29]),
        .s(fa_s0_c67_n382_s),
        .c_out(fa_s0_c67_n382_c)
    );

    fa fa_s0_c68_n383 (
        .a(stage0_col68[0]),
        .b(stage0_col68[1]),
        .c_in(stage0_col68[2]),
        .s(fa_s0_c68_n383_s),
        .c_out(fa_s0_c68_n383_c)
    );

    fa fa_s0_c68_n384 (
        .a(stage0_col68[3]),
        .b(stage0_col68[4]),
        .c_in(stage0_col68[5]),
        .s(fa_s0_c68_n384_s),
        .c_out(fa_s0_c68_n384_c)
    );

    fa fa_s0_c68_n385 (
        .a(stage0_col68[6]),
        .b(stage0_col68[7]),
        .c_in(stage0_col68[8]),
        .s(fa_s0_c68_n385_s),
        .c_out(fa_s0_c68_n385_c)
    );

    fa fa_s0_c68_n386 (
        .a(stage0_col68[9]),
        .b(stage0_col68[10]),
        .c_in(stage0_col68[11]),
        .s(fa_s0_c68_n386_s),
        .c_out(fa_s0_c68_n386_c)
    );

    fa fa_s0_c68_n387 (
        .a(stage0_col68[12]),
        .b(stage0_col68[13]),
        .c_in(stage0_col68[14]),
        .s(fa_s0_c68_n387_s),
        .c_out(fa_s0_c68_n387_c)
    );

    fa fa_s0_c68_n388 (
        .a(stage0_col68[15]),
        .b(stage0_col68[16]),
        .c_in(stage0_col68[17]),
        .s(fa_s0_c68_n388_s),
        .c_out(fa_s0_c68_n388_c)
    );

    fa fa_s0_c68_n389 (
        .a(stage0_col68[18]),
        .b(stage0_col68[19]),
        .c_in(stage0_col68[20]),
        .s(fa_s0_c68_n389_s),
        .c_out(fa_s0_c68_n389_c)
    );

    fa fa_s0_c68_n390 (
        .a(stage0_col68[21]),
        .b(stage0_col68[22]),
        .c_in(stage0_col68[23]),
        .s(fa_s0_c68_n390_s),
        .c_out(fa_s0_c68_n390_c)
    );

    fa fa_s0_c68_n391 (
        .a(stage0_col68[24]),
        .b(stage0_col68[25]),
        .c_in(stage0_col68[26]),
        .s(fa_s0_c68_n391_s),
        .c_out(fa_s0_c68_n391_c)
    );

    fa fa_s0_c68_n392 (
        .a(stage0_col68[27]),
        .b(stage0_col68[28]),
        .c_in(stage0_col68[29]),
        .s(fa_s0_c68_n392_s),
        .c_out(fa_s0_c68_n392_c)
    );

    fa fa_s0_c68_n393 (
        .a(stage0_col68[30]),
        .b(stage0_col68[31]),
        .c_in(stage0_col68[32]),
        .s(fa_s0_c68_n393_s),
        .c_out(fa_s0_c68_n393_c)
    );

    fa fa_s0_c69_n394 (
        .a(stage0_col69[0]),
        .b(stage0_col69[1]),
        .c_in(stage0_col69[2]),
        .s(fa_s0_c69_n394_s),
        .c_out(fa_s0_c69_n394_c)
    );

    fa fa_s0_c69_n395 (
        .a(stage0_col69[3]),
        .b(stage0_col69[4]),
        .c_in(stage0_col69[5]),
        .s(fa_s0_c69_n395_s),
        .c_out(fa_s0_c69_n395_c)
    );

    fa fa_s0_c69_n396 (
        .a(stage0_col69[6]),
        .b(stage0_col69[7]),
        .c_in(stage0_col69[8]),
        .s(fa_s0_c69_n396_s),
        .c_out(fa_s0_c69_n396_c)
    );

    fa fa_s0_c69_n397 (
        .a(stage0_col69[9]),
        .b(stage0_col69[10]),
        .c_in(stage0_col69[11]),
        .s(fa_s0_c69_n397_s),
        .c_out(fa_s0_c69_n397_c)
    );

    fa fa_s0_c69_n398 (
        .a(stage0_col69[12]),
        .b(stage0_col69[13]),
        .c_in(stage0_col69[14]),
        .s(fa_s0_c69_n398_s),
        .c_out(fa_s0_c69_n398_c)
    );

    fa fa_s0_c69_n399 (
        .a(stage0_col69[15]),
        .b(stage0_col69[16]),
        .c_in(stage0_col69[17]),
        .s(fa_s0_c69_n399_s),
        .c_out(fa_s0_c69_n399_c)
    );

    fa fa_s0_c69_n400 (
        .a(stage0_col69[18]),
        .b(stage0_col69[19]),
        .c_in(stage0_col69[20]),
        .s(fa_s0_c69_n400_s),
        .c_out(fa_s0_c69_n400_c)
    );

    fa fa_s0_c69_n401 (
        .a(stage0_col69[21]),
        .b(stage0_col69[22]),
        .c_in(stage0_col69[23]),
        .s(fa_s0_c69_n401_s),
        .c_out(fa_s0_c69_n401_c)
    );

    fa fa_s0_c69_n402 (
        .a(stage0_col69[24]),
        .b(stage0_col69[25]),
        .c_in(stage0_col69[26]),
        .s(fa_s0_c69_n402_s),
        .c_out(fa_s0_c69_n402_c)
    );

    fa fa_s0_c69_n403 (
        .a(stage0_col69[27]),
        .b(stage0_col69[28]),
        .c_in(stage0_col69[29]),
        .s(fa_s0_c69_n403_s),
        .c_out(fa_s0_c69_n403_c)
    );

    fa fa_s0_c70_n404 (
        .a(stage0_col70[0]),
        .b(stage0_col70[1]),
        .c_in(stage0_col70[2]),
        .s(fa_s0_c70_n404_s),
        .c_out(fa_s0_c70_n404_c)
    );

    fa fa_s0_c70_n405 (
        .a(stage0_col70[3]),
        .b(stage0_col70[4]),
        .c_in(stage0_col70[5]),
        .s(fa_s0_c70_n405_s),
        .c_out(fa_s0_c70_n405_c)
    );

    fa fa_s0_c70_n406 (
        .a(stage0_col70[6]),
        .b(stage0_col70[7]),
        .c_in(stage0_col70[8]),
        .s(fa_s0_c70_n406_s),
        .c_out(fa_s0_c70_n406_c)
    );

    fa fa_s0_c70_n407 (
        .a(stage0_col70[9]),
        .b(stage0_col70[10]),
        .c_in(stage0_col70[11]),
        .s(fa_s0_c70_n407_s),
        .c_out(fa_s0_c70_n407_c)
    );

    fa fa_s0_c70_n408 (
        .a(stage0_col70[12]),
        .b(stage0_col70[13]),
        .c_in(stage0_col70[14]),
        .s(fa_s0_c70_n408_s),
        .c_out(fa_s0_c70_n408_c)
    );

    fa fa_s0_c70_n409 (
        .a(stage0_col70[15]),
        .b(stage0_col70[16]),
        .c_in(stage0_col70[17]),
        .s(fa_s0_c70_n409_s),
        .c_out(fa_s0_c70_n409_c)
    );

    fa fa_s0_c70_n410 (
        .a(stage0_col70[18]),
        .b(stage0_col70[19]),
        .c_in(stage0_col70[20]),
        .s(fa_s0_c70_n410_s),
        .c_out(fa_s0_c70_n410_c)
    );

    fa fa_s0_c70_n411 (
        .a(stage0_col70[21]),
        .b(stage0_col70[22]),
        .c_in(stage0_col70[23]),
        .s(fa_s0_c70_n411_s),
        .c_out(fa_s0_c70_n411_c)
    );

    fa fa_s0_c70_n412 (
        .a(stage0_col70[24]),
        .b(stage0_col70[25]),
        .c_in(stage0_col70[26]),
        .s(fa_s0_c70_n412_s),
        .c_out(fa_s0_c70_n412_c)
    );

    fa fa_s0_c70_n413 (
        .a(stage0_col70[27]),
        .b(stage0_col70[28]),
        .c_in(stage0_col70[29]),
        .s(fa_s0_c70_n413_s),
        .c_out(fa_s0_c70_n413_c)
    );

    fa fa_s0_c70_n414 (
        .a(stage0_col70[30]),
        .b(stage0_col70[31]),
        .c_in(stage0_col70[32]),
        .s(fa_s0_c70_n414_s),
        .c_out(fa_s0_c70_n414_c)
    );

    fa fa_s0_c71_n415 (
        .a(stage0_col71[0]),
        .b(stage0_col71[1]),
        .c_in(stage0_col71[2]),
        .s(fa_s0_c71_n415_s),
        .c_out(fa_s0_c71_n415_c)
    );

    fa fa_s0_c71_n416 (
        .a(stage0_col71[3]),
        .b(stage0_col71[4]),
        .c_in(stage0_col71[5]),
        .s(fa_s0_c71_n416_s),
        .c_out(fa_s0_c71_n416_c)
    );

    fa fa_s0_c71_n417 (
        .a(stage0_col71[6]),
        .b(stage0_col71[7]),
        .c_in(stage0_col71[8]),
        .s(fa_s0_c71_n417_s),
        .c_out(fa_s0_c71_n417_c)
    );

    fa fa_s0_c71_n418 (
        .a(stage0_col71[9]),
        .b(stage0_col71[10]),
        .c_in(stage0_col71[11]),
        .s(fa_s0_c71_n418_s),
        .c_out(fa_s0_c71_n418_c)
    );

    fa fa_s0_c71_n419 (
        .a(stage0_col71[12]),
        .b(stage0_col71[13]),
        .c_in(stage0_col71[14]),
        .s(fa_s0_c71_n419_s),
        .c_out(fa_s0_c71_n419_c)
    );

    fa fa_s0_c71_n420 (
        .a(stage0_col71[15]),
        .b(stage0_col71[16]),
        .c_in(stage0_col71[17]),
        .s(fa_s0_c71_n420_s),
        .c_out(fa_s0_c71_n420_c)
    );

    fa fa_s0_c71_n421 (
        .a(stage0_col71[18]),
        .b(stage0_col71[19]),
        .c_in(stage0_col71[20]),
        .s(fa_s0_c71_n421_s),
        .c_out(fa_s0_c71_n421_c)
    );

    fa fa_s0_c71_n422 (
        .a(stage0_col71[21]),
        .b(stage0_col71[22]),
        .c_in(stage0_col71[23]),
        .s(fa_s0_c71_n422_s),
        .c_out(fa_s0_c71_n422_c)
    );

    fa fa_s0_c71_n423 (
        .a(stage0_col71[24]),
        .b(stage0_col71[25]),
        .c_in(stage0_col71[26]),
        .s(fa_s0_c71_n423_s),
        .c_out(fa_s0_c71_n423_c)
    );

    fa fa_s0_c71_n424 (
        .a(stage0_col71[27]),
        .b(stage0_col71[28]),
        .c_in(stage0_col71[29]),
        .s(fa_s0_c71_n424_s),
        .c_out(fa_s0_c71_n424_c)
    );

    fa fa_s0_c72_n425 (
        .a(stage0_col72[0]),
        .b(stage0_col72[1]),
        .c_in(stage0_col72[2]),
        .s(fa_s0_c72_n425_s),
        .c_out(fa_s0_c72_n425_c)
    );

    fa fa_s0_c72_n426 (
        .a(stage0_col72[3]),
        .b(stage0_col72[4]),
        .c_in(stage0_col72[5]),
        .s(fa_s0_c72_n426_s),
        .c_out(fa_s0_c72_n426_c)
    );

    fa fa_s0_c72_n427 (
        .a(stage0_col72[6]),
        .b(stage0_col72[7]),
        .c_in(stage0_col72[8]),
        .s(fa_s0_c72_n427_s),
        .c_out(fa_s0_c72_n427_c)
    );

    fa fa_s0_c72_n428 (
        .a(stage0_col72[9]),
        .b(stage0_col72[10]),
        .c_in(stage0_col72[11]),
        .s(fa_s0_c72_n428_s),
        .c_out(fa_s0_c72_n428_c)
    );

    fa fa_s0_c72_n429 (
        .a(stage0_col72[12]),
        .b(stage0_col72[13]),
        .c_in(stage0_col72[14]),
        .s(fa_s0_c72_n429_s),
        .c_out(fa_s0_c72_n429_c)
    );

    fa fa_s0_c72_n430 (
        .a(stage0_col72[15]),
        .b(stage0_col72[16]),
        .c_in(stage0_col72[17]),
        .s(fa_s0_c72_n430_s),
        .c_out(fa_s0_c72_n430_c)
    );

    fa fa_s0_c72_n431 (
        .a(stage0_col72[18]),
        .b(stage0_col72[19]),
        .c_in(stage0_col72[20]),
        .s(fa_s0_c72_n431_s),
        .c_out(fa_s0_c72_n431_c)
    );

    fa fa_s0_c72_n432 (
        .a(stage0_col72[21]),
        .b(stage0_col72[22]),
        .c_in(stage0_col72[23]),
        .s(fa_s0_c72_n432_s),
        .c_out(fa_s0_c72_n432_c)
    );

    fa fa_s0_c72_n433 (
        .a(stage0_col72[24]),
        .b(stage0_col72[25]),
        .c_in(stage0_col72[26]),
        .s(fa_s0_c72_n433_s),
        .c_out(fa_s0_c72_n433_c)
    );

    fa fa_s0_c72_n434 (
        .a(stage0_col72[27]),
        .b(stage0_col72[28]),
        .c_in(stage0_col72[29]),
        .s(fa_s0_c72_n434_s),
        .c_out(fa_s0_c72_n434_c)
    );

    fa fa_s0_c72_n435 (
        .a(stage0_col72[30]),
        .b(stage0_col72[31]),
        .c_in(stage0_col72[32]),
        .s(fa_s0_c72_n435_s),
        .c_out(fa_s0_c72_n435_c)
    );

    fa fa_s0_c73_n436 (
        .a(stage0_col73[0]),
        .b(stage0_col73[1]),
        .c_in(stage0_col73[2]),
        .s(fa_s0_c73_n436_s),
        .c_out(fa_s0_c73_n436_c)
    );

    fa fa_s0_c73_n437 (
        .a(stage0_col73[3]),
        .b(stage0_col73[4]),
        .c_in(stage0_col73[5]),
        .s(fa_s0_c73_n437_s),
        .c_out(fa_s0_c73_n437_c)
    );

    fa fa_s0_c73_n438 (
        .a(stage0_col73[6]),
        .b(stage0_col73[7]),
        .c_in(stage0_col73[8]),
        .s(fa_s0_c73_n438_s),
        .c_out(fa_s0_c73_n438_c)
    );

    fa fa_s0_c73_n439 (
        .a(stage0_col73[9]),
        .b(stage0_col73[10]),
        .c_in(stage0_col73[11]),
        .s(fa_s0_c73_n439_s),
        .c_out(fa_s0_c73_n439_c)
    );

    fa fa_s0_c73_n440 (
        .a(stage0_col73[12]),
        .b(stage0_col73[13]),
        .c_in(stage0_col73[14]),
        .s(fa_s0_c73_n440_s),
        .c_out(fa_s0_c73_n440_c)
    );

    fa fa_s0_c73_n441 (
        .a(stage0_col73[15]),
        .b(stage0_col73[16]),
        .c_in(stage0_col73[17]),
        .s(fa_s0_c73_n441_s),
        .c_out(fa_s0_c73_n441_c)
    );

    fa fa_s0_c73_n442 (
        .a(stage0_col73[18]),
        .b(stage0_col73[19]),
        .c_in(stage0_col73[20]),
        .s(fa_s0_c73_n442_s),
        .c_out(fa_s0_c73_n442_c)
    );

    fa fa_s0_c73_n443 (
        .a(stage0_col73[21]),
        .b(stage0_col73[22]),
        .c_in(stage0_col73[23]),
        .s(fa_s0_c73_n443_s),
        .c_out(fa_s0_c73_n443_c)
    );

    fa fa_s0_c73_n444 (
        .a(stage0_col73[24]),
        .b(stage0_col73[25]),
        .c_in(stage0_col73[26]),
        .s(fa_s0_c73_n444_s),
        .c_out(fa_s0_c73_n444_c)
    );

    fa fa_s0_c73_n445 (
        .a(stage0_col73[27]),
        .b(stage0_col73[28]),
        .c_in(stage0_col73[29]),
        .s(fa_s0_c73_n445_s),
        .c_out(fa_s0_c73_n445_c)
    );

    fa fa_s0_c74_n446 (
        .a(stage0_col74[0]),
        .b(stage0_col74[1]),
        .c_in(stage0_col74[2]),
        .s(fa_s0_c74_n446_s),
        .c_out(fa_s0_c74_n446_c)
    );

    fa fa_s0_c74_n447 (
        .a(stage0_col74[3]),
        .b(stage0_col74[4]),
        .c_in(stage0_col74[5]),
        .s(fa_s0_c74_n447_s),
        .c_out(fa_s0_c74_n447_c)
    );

    fa fa_s0_c74_n448 (
        .a(stage0_col74[6]),
        .b(stage0_col74[7]),
        .c_in(stage0_col74[8]),
        .s(fa_s0_c74_n448_s),
        .c_out(fa_s0_c74_n448_c)
    );

    fa fa_s0_c74_n449 (
        .a(stage0_col74[9]),
        .b(stage0_col74[10]),
        .c_in(stage0_col74[11]),
        .s(fa_s0_c74_n449_s),
        .c_out(fa_s0_c74_n449_c)
    );

    fa fa_s0_c74_n450 (
        .a(stage0_col74[12]),
        .b(stage0_col74[13]),
        .c_in(stage0_col74[14]),
        .s(fa_s0_c74_n450_s),
        .c_out(fa_s0_c74_n450_c)
    );

    fa fa_s0_c74_n451 (
        .a(stage0_col74[15]),
        .b(stage0_col74[16]),
        .c_in(stage0_col74[17]),
        .s(fa_s0_c74_n451_s),
        .c_out(fa_s0_c74_n451_c)
    );

    fa fa_s0_c74_n452 (
        .a(stage0_col74[18]),
        .b(stage0_col74[19]),
        .c_in(stage0_col74[20]),
        .s(fa_s0_c74_n452_s),
        .c_out(fa_s0_c74_n452_c)
    );

    fa fa_s0_c74_n453 (
        .a(stage0_col74[21]),
        .b(stage0_col74[22]),
        .c_in(stage0_col74[23]),
        .s(fa_s0_c74_n453_s),
        .c_out(fa_s0_c74_n453_c)
    );

    fa fa_s0_c74_n454 (
        .a(stage0_col74[24]),
        .b(stage0_col74[25]),
        .c_in(stage0_col74[26]),
        .s(fa_s0_c74_n454_s),
        .c_out(fa_s0_c74_n454_c)
    );

    fa fa_s0_c74_n455 (
        .a(stage0_col74[27]),
        .b(stage0_col74[28]),
        .c_in(stage0_col74[29]),
        .s(fa_s0_c74_n455_s),
        .c_out(fa_s0_c74_n455_c)
    );

    fa fa_s0_c74_n456 (
        .a(stage0_col74[30]),
        .b(stage0_col74[31]),
        .c_in(stage0_col74[32]),
        .s(fa_s0_c74_n456_s),
        .c_out(fa_s0_c74_n456_c)
    );

    fa fa_s0_c75_n457 (
        .a(stage0_col75[0]),
        .b(stage0_col75[1]),
        .c_in(stage0_col75[2]),
        .s(fa_s0_c75_n457_s),
        .c_out(fa_s0_c75_n457_c)
    );

    fa fa_s0_c75_n458 (
        .a(stage0_col75[3]),
        .b(stage0_col75[4]),
        .c_in(stage0_col75[5]),
        .s(fa_s0_c75_n458_s),
        .c_out(fa_s0_c75_n458_c)
    );

    fa fa_s0_c75_n459 (
        .a(stage0_col75[6]),
        .b(stage0_col75[7]),
        .c_in(stage0_col75[8]),
        .s(fa_s0_c75_n459_s),
        .c_out(fa_s0_c75_n459_c)
    );

    fa fa_s0_c75_n460 (
        .a(stage0_col75[9]),
        .b(stage0_col75[10]),
        .c_in(stage0_col75[11]),
        .s(fa_s0_c75_n460_s),
        .c_out(fa_s0_c75_n460_c)
    );

    fa fa_s0_c75_n461 (
        .a(stage0_col75[12]),
        .b(stage0_col75[13]),
        .c_in(stage0_col75[14]),
        .s(fa_s0_c75_n461_s),
        .c_out(fa_s0_c75_n461_c)
    );

    fa fa_s0_c75_n462 (
        .a(stage0_col75[15]),
        .b(stage0_col75[16]),
        .c_in(stage0_col75[17]),
        .s(fa_s0_c75_n462_s),
        .c_out(fa_s0_c75_n462_c)
    );

    fa fa_s0_c75_n463 (
        .a(stage0_col75[18]),
        .b(stage0_col75[19]),
        .c_in(stage0_col75[20]),
        .s(fa_s0_c75_n463_s),
        .c_out(fa_s0_c75_n463_c)
    );

    fa fa_s0_c75_n464 (
        .a(stage0_col75[21]),
        .b(stage0_col75[22]),
        .c_in(stage0_col75[23]),
        .s(fa_s0_c75_n464_s),
        .c_out(fa_s0_c75_n464_c)
    );

    fa fa_s0_c75_n465 (
        .a(stage0_col75[24]),
        .b(stage0_col75[25]),
        .c_in(stage0_col75[26]),
        .s(fa_s0_c75_n465_s),
        .c_out(fa_s0_c75_n465_c)
    );

    fa fa_s0_c75_n466 (
        .a(stage0_col75[27]),
        .b(stage0_col75[28]),
        .c_in(stage0_col75[29]),
        .s(fa_s0_c75_n466_s),
        .c_out(fa_s0_c75_n466_c)
    );

    fa fa_s0_c76_n467 (
        .a(stage0_col76[0]),
        .b(stage0_col76[1]),
        .c_in(stage0_col76[2]),
        .s(fa_s0_c76_n467_s),
        .c_out(fa_s0_c76_n467_c)
    );

    fa fa_s0_c76_n468 (
        .a(stage0_col76[3]),
        .b(stage0_col76[4]),
        .c_in(stage0_col76[5]),
        .s(fa_s0_c76_n468_s),
        .c_out(fa_s0_c76_n468_c)
    );

    fa fa_s0_c76_n469 (
        .a(stage0_col76[6]),
        .b(stage0_col76[7]),
        .c_in(stage0_col76[8]),
        .s(fa_s0_c76_n469_s),
        .c_out(fa_s0_c76_n469_c)
    );

    fa fa_s0_c76_n470 (
        .a(stage0_col76[9]),
        .b(stage0_col76[10]),
        .c_in(stage0_col76[11]),
        .s(fa_s0_c76_n470_s),
        .c_out(fa_s0_c76_n470_c)
    );

    fa fa_s0_c76_n471 (
        .a(stage0_col76[12]),
        .b(stage0_col76[13]),
        .c_in(stage0_col76[14]),
        .s(fa_s0_c76_n471_s),
        .c_out(fa_s0_c76_n471_c)
    );

    fa fa_s0_c76_n472 (
        .a(stage0_col76[15]),
        .b(stage0_col76[16]),
        .c_in(stage0_col76[17]),
        .s(fa_s0_c76_n472_s),
        .c_out(fa_s0_c76_n472_c)
    );

    fa fa_s0_c76_n473 (
        .a(stage0_col76[18]),
        .b(stage0_col76[19]),
        .c_in(stage0_col76[20]),
        .s(fa_s0_c76_n473_s),
        .c_out(fa_s0_c76_n473_c)
    );

    fa fa_s0_c76_n474 (
        .a(stage0_col76[21]),
        .b(stage0_col76[22]),
        .c_in(stage0_col76[23]),
        .s(fa_s0_c76_n474_s),
        .c_out(fa_s0_c76_n474_c)
    );

    fa fa_s0_c76_n475 (
        .a(stage0_col76[24]),
        .b(stage0_col76[25]),
        .c_in(stage0_col76[26]),
        .s(fa_s0_c76_n475_s),
        .c_out(fa_s0_c76_n475_c)
    );

    fa fa_s0_c76_n476 (
        .a(stage0_col76[27]),
        .b(stage0_col76[28]),
        .c_in(stage0_col76[29]),
        .s(fa_s0_c76_n476_s),
        .c_out(fa_s0_c76_n476_c)
    );

    fa fa_s0_c76_n477 (
        .a(stage0_col76[30]),
        .b(stage0_col76[31]),
        .c_in(stage0_col76[32]),
        .s(fa_s0_c76_n477_s),
        .c_out(fa_s0_c76_n477_c)
    );

    fa fa_s0_c77_n478 (
        .a(stage0_col77[0]),
        .b(stage0_col77[1]),
        .c_in(stage0_col77[2]),
        .s(fa_s0_c77_n478_s),
        .c_out(fa_s0_c77_n478_c)
    );

    fa fa_s0_c77_n479 (
        .a(stage0_col77[3]),
        .b(stage0_col77[4]),
        .c_in(stage0_col77[5]),
        .s(fa_s0_c77_n479_s),
        .c_out(fa_s0_c77_n479_c)
    );

    fa fa_s0_c77_n480 (
        .a(stage0_col77[6]),
        .b(stage0_col77[7]),
        .c_in(stage0_col77[8]),
        .s(fa_s0_c77_n480_s),
        .c_out(fa_s0_c77_n480_c)
    );

    fa fa_s0_c77_n481 (
        .a(stage0_col77[9]),
        .b(stage0_col77[10]),
        .c_in(stage0_col77[11]),
        .s(fa_s0_c77_n481_s),
        .c_out(fa_s0_c77_n481_c)
    );

    fa fa_s0_c77_n482 (
        .a(stage0_col77[12]),
        .b(stage0_col77[13]),
        .c_in(stage0_col77[14]),
        .s(fa_s0_c77_n482_s),
        .c_out(fa_s0_c77_n482_c)
    );

    fa fa_s0_c77_n483 (
        .a(stage0_col77[15]),
        .b(stage0_col77[16]),
        .c_in(stage0_col77[17]),
        .s(fa_s0_c77_n483_s),
        .c_out(fa_s0_c77_n483_c)
    );

    fa fa_s0_c77_n484 (
        .a(stage0_col77[18]),
        .b(stage0_col77[19]),
        .c_in(stage0_col77[20]),
        .s(fa_s0_c77_n484_s),
        .c_out(fa_s0_c77_n484_c)
    );

    fa fa_s0_c77_n485 (
        .a(stage0_col77[21]),
        .b(stage0_col77[22]),
        .c_in(stage0_col77[23]),
        .s(fa_s0_c77_n485_s),
        .c_out(fa_s0_c77_n485_c)
    );

    fa fa_s0_c77_n486 (
        .a(stage0_col77[24]),
        .b(stage0_col77[25]),
        .c_in(stage0_col77[26]),
        .s(fa_s0_c77_n486_s),
        .c_out(fa_s0_c77_n486_c)
    );

    fa fa_s0_c77_n487 (
        .a(stage0_col77[27]),
        .b(stage0_col77[28]),
        .c_in(stage0_col77[29]),
        .s(fa_s0_c77_n487_s),
        .c_out(fa_s0_c77_n487_c)
    );

    fa fa_s0_c78_n488 (
        .a(stage0_col78[0]),
        .b(stage0_col78[1]),
        .c_in(stage0_col78[2]),
        .s(fa_s0_c78_n488_s),
        .c_out(fa_s0_c78_n488_c)
    );

    fa fa_s0_c78_n489 (
        .a(stage0_col78[3]),
        .b(stage0_col78[4]),
        .c_in(stage0_col78[5]),
        .s(fa_s0_c78_n489_s),
        .c_out(fa_s0_c78_n489_c)
    );

    fa fa_s0_c78_n490 (
        .a(stage0_col78[6]),
        .b(stage0_col78[7]),
        .c_in(stage0_col78[8]),
        .s(fa_s0_c78_n490_s),
        .c_out(fa_s0_c78_n490_c)
    );

    fa fa_s0_c78_n491 (
        .a(stage0_col78[9]),
        .b(stage0_col78[10]),
        .c_in(stage0_col78[11]),
        .s(fa_s0_c78_n491_s),
        .c_out(fa_s0_c78_n491_c)
    );

    fa fa_s0_c78_n492 (
        .a(stage0_col78[12]),
        .b(stage0_col78[13]),
        .c_in(stage0_col78[14]),
        .s(fa_s0_c78_n492_s),
        .c_out(fa_s0_c78_n492_c)
    );

    fa fa_s0_c78_n493 (
        .a(stage0_col78[15]),
        .b(stage0_col78[16]),
        .c_in(stage0_col78[17]),
        .s(fa_s0_c78_n493_s),
        .c_out(fa_s0_c78_n493_c)
    );

    fa fa_s0_c78_n494 (
        .a(stage0_col78[18]),
        .b(stage0_col78[19]),
        .c_in(stage0_col78[20]),
        .s(fa_s0_c78_n494_s),
        .c_out(fa_s0_c78_n494_c)
    );

    fa fa_s0_c78_n495 (
        .a(stage0_col78[21]),
        .b(stage0_col78[22]),
        .c_in(stage0_col78[23]),
        .s(fa_s0_c78_n495_s),
        .c_out(fa_s0_c78_n495_c)
    );

    fa fa_s0_c78_n496 (
        .a(stage0_col78[24]),
        .b(stage0_col78[25]),
        .c_in(stage0_col78[26]),
        .s(fa_s0_c78_n496_s),
        .c_out(fa_s0_c78_n496_c)
    );

    fa fa_s0_c78_n497 (
        .a(stage0_col78[27]),
        .b(stage0_col78[28]),
        .c_in(stage0_col78[29]),
        .s(fa_s0_c78_n497_s),
        .c_out(fa_s0_c78_n497_c)
    );

    fa fa_s0_c78_n498 (
        .a(stage0_col78[30]),
        .b(stage0_col78[31]),
        .c_in(stage0_col78[32]),
        .s(fa_s0_c78_n498_s),
        .c_out(fa_s0_c78_n498_c)
    );

    fa fa_s0_c79_n499 (
        .a(stage0_col79[0]),
        .b(stage0_col79[1]),
        .c_in(stage0_col79[2]),
        .s(fa_s0_c79_n499_s),
        .c_out(fa_s0_c79_n499_c)
    );

    fa fa_s0_c79_n500 (
        .a(stage0_col79[3]),
        .b(stage0_col79[4]),
        .c_in(stage0_col79[5]),
        .s(fa_s0_c79_n500_s),
        .c_out(fa_s0_c79_n500_c)
    );

    fa fa_s0_c79_n501 (
        .a(stage0_col79[6]),
        .b(stage0_col79[7]),
        .c_in(stage0_col79[8]),
        .s(fa_s0_c79_n501_s),
        .c_out(fa_s0_c79_n501_c)
    );

    fa fa_s0_c79_n502 (
        .a(stage0_col79[9]),
        .b(stage0_col79[10]),
        .c_in(stage0_col79[11]),
        .s(fa_s0_c79_n502_s),
        .c_out(fa_s0_c79_n502_c)
    );

    fa fa_s0_c79_n503 (
        .a(stage0_col79[12]),
        .b(stage0_col79[13]),
        .c_in(stage0_col79[14]),
        .s(fa_s0_c79_n503_s),
        .c_out(fa_s0_c79_n503_c)
    );

    fa fa_s0_c79_n504 (
        .a(stage0_col79[15]),
        .b(stage0_col79[16]),
        .c_in(stage0_col79[17]),
        .s(fa_s0_c79_n504_s),
        .c_out(fa_s0_c79_n504_c)
    );

    fa fa_s0_c79_n505 (
        .a(stage0_col79[18]),
        .b(stage0_col79[19]),
        .c_in(stage0_col79[20]),
        .s(fa_s0_c79_n505_s),
        .c_out(fa_s0_c79_n505_c)
    );

    fa fa_s0_c79_n506 (
        .a(stage0_col79[21]),
        .b(stage0_col79[22]),
        .c_in(stage0_col79[23]),
        .s(fa_s0_c79_n506_s),
        .c_out(fa_s0_c79_n506_c)
    );

    fa fa_s0_c79_n507 (
        .a(stage0_col79[24]),
        .b(stage0_col79[25]),
        .c_in(stage0_col79[26]),
        .s(fa_s0_c79_n507_s),
        .c_out(fa_s0_c79_n507_c)
    );

    fa fa_s0_c79_n508 (
        .a(stage0_col79[27]),
        .b(stage0_col79[28]),
        .c_in(stage0_col79[29]),
        .s(fa_s0_c79_n508_s),
        .c_out(fa_s0_c79_n508_c)
    );

    fa fa_s0_c80_n509 (
        .a(stage0_col80[0]),
        .b(stage0_col80[1]),
        .c_in(stage0_col80[2]),
        .s(fa_s0_c80_n509_s),
        .c_out(fa_s0_c80_n509_c)
    );

    fa fa_s0_c80_n510 (
        .a(stage0_col80[3]),
        .b(stage0_col80[4]),
        .c_in(stage0_col80[5]),
        .s(fa_s0_c80_n510_s),
        .c_out(fa_s0_c80_n510_c)
    );

    fa fa_s0_c80_n511 (
        .a(stage0_col80[6]),
        .b(stage0_col80[7]),
        .c_in(stage0_col80[8]),
        .s(fa_s0_c80_n511_s),
        .c_out(fa_s0_c80_n511_c)
    );

    fa fa_s0_c80_n512 (
        .a(stage0_col80[9]),
        .b(stage0_col80[10]),
        .c_in(stage0_col80[11]),
        .s(fa_s0_c80_n512_s),
        .c_out(fa_s0_c80_n512_c)
    );

    fa fa_s0_c80_n513 (
        .a(stage0_col80[12]),
        .b(stage0_col80[13]),
        .c_in(stage0_col80[14]),
        .s(fa_s0_c80_n513_s),
        .c_out(fa_s0_c80_n513_c)
    );

    fa fa_s0_c80_n514 (
        .a(stage0_col80[15]),
        .b(stage0_col80[16]),
        .c_in(stage0_col80[17]),
        .s(fa_s0_c80_n514_s),
        .c_out(fa_s0_c80_n514_c)
    );

    fa fa_s0_c80_n515 (
        .a(stage0_col80[18]),
        .b(stage0_col80[19]),
        .c_in(stage0_col80[20]),
        .s(fa_s0_c80_n515_s),
        .c_out(fa_s0_c80_n515_c)
    );

    fa fa_s0_c80_n516 (
        .a(stage0_col80[21]),
        .b(stage0_col80[22]),
        .c_in(stage0_col80[23]),
        .s(fa_s0_c80_n516_s),
        .c_out(fa_s0_c80_n516_c)
    );

    fa fa_s0_c80_n517 (
        .a(stage0_col80[24]),
        .b(stage0_col80[25]),
        .c_in(stage0_col80[26]),
        .s(fa_s0_c80_n517_s),
        .c_out(fa_s0_c80_n517_c)
    );

    fa fa_s0_c80_n518 (
        .a(stage0_col80[27]),
        .b(stage0_col80[28]),
        .c_in(stage0_col80[29]),
        .s(fa_s0_c80_n518_s),
        .c_out(fa_s0_c80_n518_c)
    );

    fa fa_s0_c80_n519 (
        .a(stage0_col80[30]),
        .b(stage0_col80[31]),
        .c_in(stage0_col80[32]),
        .s(fa_s0_c80_n519_s),
        .c_out(fa_s0_c80_n519_c)
    );

    fa fa_s0_c81_n520 (
        .a(stage0_col81[0]),
        .b(stage0_col81[1]),
        .c_in(stage0_col81[2]),
        .s(fa_s0_c81_n520_s),
        .c_out(fa_s0_c81_n520_c)
    );

    fa fa_s0_c81_n521 (
        .a(stage0_col81[3]),
        .b(stage0_col81[4]),
        .c_in(stage0_col81[5]),
        .s(fa_s0_c81_n521_s),
        .c_out(fa_s0_c81_n521_c)
    );

    fa fa_s0_c81_n522 (
        .a(stage0_col81[6]),
        .b(stage0_col81[7]),
        .c_in(stage0_col81[8]),
        .s(fa_s0_c81_n522_s),
        .c_out(fa_s0_c81_n522_c)
    );

    fa fa_s0_c81_n523 (
        .a(stage0_col81[9]),
        .b(stage0_col81[10]),
        .c_in(stage0_col81[11]),
        .s(fa_s0_c81_n523_s),
        .c_out(fa_s0_c81_n523_c)
    );

    fa fa_s0_c81_n524 (
        .a(stage0_col81[12]),
        .b(stage0_col81[13]),
        .c_in(stage0_col81[14]),
        .s(fa_s0_c81_n524_s),
        .c_out(fa_s0_c81_n524_c)
    );

    fa fa_s0_c81_n525 (
        .a(stage0_col81[15]),
        .b(stage0_col81[16]),
        .c_in(stage0_col81[17]),
        .s(fa_s0_c81_n525_s),
        .c_out(fa_s0_c81_n525_c)
    );

    fa fa_s0_c81_n526 (
        .a(stage0_col81[18]),
        .b(stage0_col81[19]),
        .c_in(stage0_col81[20]),
        .s(fa_s0_c81_n526_s),
        .c_out(fa_s0_c81_n526_c)
    );

    fa fa_s0_c81_n527 (
        .a(stage0_col81[21]),
        .b(stage0_col81[22]),
        .c_in(stage0_col81[23]),
        .s(fa_s0_c81_n527_s),
        .c_out(fa_s0_c81_n527_c)
    );

    fa fa_s0_c81_n528 (
        .a(stage0_col81[24]),
        .b(stage0_col81[25]),
        .c_in(stage0_col81[26]),
        .s(fa_s0_c81_n528_s),
        .c_out(fa_s0_c81_n528_c)
    );

    fa fa_s0_c81_n529 (
        .a(stage0_col81[27]),
        .b(stage0_col81[28]),
        .c_in(stage0_col81[29]),
        .s(fa_s0_c81_n529_s),
        .c_out(fa_s0_c81_n529_c)
    );

    fa fa_s0_c82_n530 (
        .a(stage0_col82[0]),
        .b(stage0_col82[1]),
        .c_in(stage0_col82[2]),
        .s(fa_s0_c82_n530_s),
        .c_out(fa_s0_c82_n530_c)
    );

    fa fa_s0_c82_n531 (
        .a(stage0_col82[3]),
        .b(stage0_col82[4]),
        .c_in(stage0_col82[5]),
        .s(fa_s0_c82_n531_s),
        .c_out(fa_s0_c82_n531_c)
    );

    fa fa_s0_c82_n532 (
        .a(stage0_col82[6]),
        .b(stage0_col82[7]),
        .c_in(stage0_col82[8]),
        .s(fa_s0_c82_n532_s),
        .c_out(fa_s0_c82_n532_c)
    );

    fa fa_s0_c82_n533 (
        .a(stage0_col82[9]),
        .b(stage0_col82[10]),
        .c_in(stage0_col82[11]),
        .s(fa_s0_c82_n533_s),
        .c_out(fa_s0_c82_n533_c)
    );

    fa fa_s0_c82_n534 (
        .a(stage0_col82[12]),
        .b(stage0_col82[13]),
        .c_in(stage0_col82[14]),
        .s(fa_s0_c82_n534_s),
        .c_out(fa_s0_c82_n534_c)
    );

    fa fa_s0_c82_n535 (
        .a(stage0_col82[15]),
        .b(stage0_col82[16]),
        .c_in(stage0_col82[17]),
        .s(fa_s0_c82_n535_s),
        .c_out(fa_s0_c82_n535_c)
    );

    fa fa_s0_c82_n536 (
        .a(stage0_col82[18]),
        .b(stage0_col82[19]),
        .c_in(stage0_col82[20]),
        .s(fa_s0_c82_n536_s),
        .c_out(fa_s0_c82_n536_c)
    );

    fa fa_s0_c82_n537 (
        .a(stage0_col82[21]),
        .b(stage0_col82[22]),
        .c_in(stage0_col82[23]),
        .s(fa_s0_c82_n537_s),
        .c_out(fa_s0_c82_n537_c)
    );

    fa fa_s0_c82_n538 (
        .a(stage0_col82[24]),
        .b(stage0_col82[25]),
        .c_in(stage0_col82[26]),
        .s(fa_s0_c82_n538_s),
        .c_out(fa_s0_c82_n538_c)
    );

    fa fa_s0_c82_n539 (
        .a(stage0_col82[27]),
        .b(stage0_col82[28]),
        .c_in(stage0_col82[29]),
        .s(fa_s0_c82_n539_s),
        .c_out(fa_s0_c82_n539_c)
    );

    fa fa_s0_c82_n540 (
        .a(stage0_col82[30]),
        .b(stage0_col82[31]),
        .c_in(stage0_col82[32]),
        .s(fa_s0_c82_n540_s),
        .c_out(fa_s0_c82_n540_c)
    );

    fa fa_s0_c83_n541 (
        .a(stage0_col83[0]),
        .b(stage0_col83[1]),
        .c_in(stage0_col83[2]),
        .s(fa_s0_c83_n541_s),
        .c_out(fa_s0_c83_n541_c)
    );

    fa fa_s0_c83_n542 (
        .a(stage0_col83[3]),
        .b(stage0_col83[4]),
        .c_in(stage0_col83[5]),
        .s(fa_s0_c83_n542_s),
        .c_out(fa_s0_c83_n542_c)
    );

    fa fa_s0_c83_n543 (
        .a(stage0_col83[6]),
        .b(stage0_col83[7]),
        .c_in(stage0_col83[8]),
        .s(fa_s0_c83_n543_s),
        .c_out(fa_s0_c83_n543_c)
    );

    fa fa_s0_c83_n544 (
        .a(stage0_col83[9]),
        .b(stage0_col83[10]),
        .c_in(stage0_col83[11]),
        .s(fa_s0_c83_n544_s),
        .c_out(fa_s0_c83_n544_c)
    );

    fa fa_s0_c83_n545 (
        .a(stage0_col83[12]),
        .b(stage0_col83[13]),
        .c_in(stage0_col83[14]),
        .s(fa_s0_c83_n545_s),
        .c_out(fa_s0_c83_n545_c)
    );

    fa fa_s0_c83_n546 (
        .a(stage0_col83[15]),
        .b(stage0_col83[16]),
        .c_in(stage0_col83[17]),
        .s(fa_s0_c83_n546_s),
        .c_out(fa_s0_c83_n546_c)
    );

    fa fa_s0_c83_n547 (
        .a(stage0_col83[18]),
        .b(stage0_col83[19]),
        .c_in(stage0_col83[20]),
        .s(fa_s0_c83_n547_s),
        .c_out(fa_s0_c83_n547_c)
    );

    fa fa_s0_c83_n548 (
        .a(stage0_col83[21]),
        .b(stage0_col83[22]),
        .c_in(stage0_col83[23]),
        .s(fa_s0_c83_n548_s),
        .c_out(fa_s0_c83_n548_c)
    );

    fa fa_s0_c83_n549 (
        .a(stage0_col83[24]),
        .b(stage0_col83[25]),
        .c_in(stage0_col83[26]),
        .s(fa_s0_c83_n549_s),
        .c_out(fa_s0_c83_n549_c)
    );

    fa fa_s0_c83_n550 (
        .a(stage0_col83[27]),
        .b(stage0_col83[28]),
        .c_in(stage0_col83[29]),
        .s(fa_s0_c83_n550_s),
        .c_out(fa_s0_c83_n550_c)
    );

    fa fa_s0_c84_n551 (
        .a(stage0_col84[0]),
        .b(stage0_col84[1]),
        .c_in(stage0_col84[2]),
        .s(fa_s0_c84_n551_s),
        .c_out(fa_s0_c84_n551_c)
    );

    fa fa_s0_c84_n552 (
        .a(stage0_col84[3]),
        .b(stage0_col84[4]),
        .c_in(stage0_col84[5]),
        .s(fa_s0_c84_n552_s),
        .c_out(fa_s0_c84_n552_c)
    );

    fa fa_s0_c84_n553 (
        .a(stage0_col84[6]),
        .b(stage0_col84[7]),
        .c_in(stage0_col84[8]),
        .s(fa_s0_c84_n553_s),
        .c_out(fa_s0_c84_n553_c)
    );

    fa fa_s0_c84_n554 (
        .a(stage0_col84[9]),
        .b(stage0_col84[10]),
        .c_in(stage0_col84[11]),
        .s(fa_s0_c84_n554_s),
        .c_out(fa_s0_c84_n554_c)
    );

    fa fa_s0_c84_n555 (
        .a(stage0_col84[12]),
        .b(stage0_col84[13]),
        .c_in(stage0_col84[14]),
        .s(fa_s0_c84_n555_s),
        .c_out(fa_s0_c84_n555_c)
    );

    fa fa_s0_c84_n556 (
        .a(stage0_col84[15]),
        .b(stage0_col84[16]),
        .c_in(stage0_col84[17]),
        .s(fa_s0_c84_n556_s),
        .c_out(fa_s0_c84_n556_c)
    );

    fa fa_s0_c84_n557 (
        .a(stage0_col84[18]),
        .b(stage0_col84[19]),
        .c_in(stage0_col84[20]),
        .s(fa_s0_c84_n557_s),
        .c_out(fa_s0_c84_n557_c)
    );

    fa fa_s0_c84_n558 (
        .a(stage0_col84[21]),
        .b(stage0_col84[22]),
        .c_in(stage0_col84[23]),
        .s(fa_s0_c84_n558_s),
        .c_out(fa_s0_c84_n558_c)
    );

    fa fa_s0_c84_n559 (
        .a(stage0_col84[24]),
        .b(stage0_col84[25]),
        .c_in(stage0_col84[26]),
        .s(fa_s0_c84_n559_s),
        .c_out(fa_s0_c84_n559_c)
    );

    fa fa_s0_c84_n560 (
        .a(stage0_col84[27]),
        .b(stage0_col84[28]),
        .c_in(stage0_col84[29]),
        .s(fa_s0_c84_n560_s),
        .c_out(fa_s0_c84_n560_c)
    );

    fa fa_s0_c84_n561 (
        .a(stage0_col84[30]),
        .b(stage0_col84[31]),
        .c_in(stage0_col84[32]),
        .s(fa_s0_c84_n561_s),
        .c_out(fa_s0_c84_n561_c)
    );

    fa fa_s0_c85_n562 (
        .a(stage0_col85[0]),
        .b(stage0_col85[1]),
        .c_in(stage0_col85[2]),
        .s(fa_s0_c85_n562_s),
        .c_out(fa_s0_c85_n562_c)
    );

    fa fa_s0_c85_n563 (
        .a(stage0_col85[3]),
        .b(stage0_col85[4]),
        .c_in(stage0_col85[5]),
        .s(fa_s0_c85_n563_s),
        .c_out(fa_s0_c85_n563_c)
    );

    fa fa_s0_c85_n564 (
        .a(stage0_col85[6]),
        .b(stage0_col85[7]),
        .c_in(stage0_col85[8]),
        .s(fa_s0_c85_n564_s),
        .c_out(fa_s0_c85_n564_c)
    );

    fa fa_s0_c85_n565 (
        .a(stage0_col85[9]),
        .b(stage0_col85[10]),
        .c_in(stage0_col85[11]),
        .s(fa_s0_c85_n565_s),
        .c_out(fa_s0_c85_n565_c)
    );

    fa fa_s0_c85_n566 (
        .a(stage0_col85[12]),
        .b(stage0_col85[13]),
        .c_in(stage0_col85[14]),
        .s(fa_s0_c85_n566_s),
        .c_out(fa_s0_c85_n566_c)
    );

    fa fa_s0_c85_n567 (
        .a(stage0_col85[15]),
        .b(stage0_col85[16]),
        .c_in(stage0_col85[17]),
        .s(fa_s0_c85_n567_s),
        .c_out(fa_s0_c85_n567_c)
    );

    fa fa_s0_c85_n568 (
        .a(stage0_col85[18]),
        .b(stage0_col85[19]),
        .c_in(stage0_col85[20]),
        .s(fa_s0_c85_n568_s),
        .c_out(fa_s0_c85_n568_c)
    );

    fa fa_s0_c85_n569 (
        .a(stage0_col85[21]),
        .b(stage0_col85[22]),
        .c_in(stage0_col85[23]),
        .s(fa_s0_c85_n569_s),
        .c_out(fa_s0_c85_n569_c)
    );

    fa fa_s0_c85_n570 (
        .a(stage0_col85[24]),
        .b(stage0_col85[25]),
        .c_in(stage0_col85[26]),
        .s(fa_s0_c85_n570_s),
        .c_out(fa_s0_c85_n570_c)
    );

    fa fa_s0_c85_n571 (
        .a(stage0_col85[27]),
        .b(stage0_col85[28]),
        .c_in(stage0_col85[29]),
        .s(fa_s0_c85_n571_s),
        .c_out(fa_s0_c85_n571_c)
    );

    fa fa_s0_c86_n572 (
        .a(stage0_col86[0]),
        .b(stage0_col86[1]),
        .c_in(stage0_col86[2]),
        .s(fa_s0_c86_n572_s),
        .c_out(fa_s0_c86_n572_c)
    );

    fa fa_s0_c86_n573 (
        .a(stage0_col86[3]),
        .b(stage0_col86[4]),
        .c_in(stage0_col86[5]),
        .s(fa_s0_c86_n573_s),
        .c_out(fa_s0_c86_n573_c)
    );

    fa fa_s0_c86_n574 (
        .a(stage0_col86[6]),
        .b(stage0_col86[7]),
        .c_in(stage0_col86[8]),
        .s(fa_s0_c86_n574_s),
        .c_out(fa_s0_c86_n574_c)
    );

    fa fa_s0_c86_n575 (
        .a(stage0_col86[9]),
        .b(stage0_col86[10]),
        .c_in(stage0_col86[11]),
        .s(fa_s0_c86_n575_s),
        .c_out(fa_s0_c86_n575_c)
    );

    fa fa_s0_c86_n576 (
        .a(stage0_col86[12]),
        .b(stage0_col86[13]),
        .c_in(stage0_col86[14]),
        .s(fa_s0_c86_n576_s),
        .c_out(fa_s0_c86_n576_c)
    );

    fa fa_s0_c86_n577 (
        .a(stage0_col86[15]),
        .b(stage0_col86[16]),
        .c_in(stage0_col86[17]),
        .s(fa_s0_c86_n577_s),
        .c_out(fa_s0_c86_n577_c)
    );

    fa fa_s0_c86_n578 (
        .a(stage0_col86[18]),
        .b(stage0_col86[19]),
        .c_in(stage0_col86[20]),
        .s(fa_s0_c86_n578_s),
        .c_out(fa_s0_c86_n578_c)
    );

    fa fa_s0_c86_n579 (
        .a(stage0_col86[21]),
        .b(stage0_col86[22]),
        .c_in(stage0_col86[23]),
        .s(fa_s0_c86_n579_s),
        .c_out(fa_s0_c86_n579_c)
    );

    fa fa_s0_c86_n580 (
        .a(stage0_col86[24]),
        .b(stage0_col86[25]),
        .c_in(stage0_col86[26]),
        .s(fa_s0_c86_n580_s),
        .c_out(fa_s0_c86_n580_c)
    );

    fa fa_s0_c86_n581 (
        .a(stage0_col86[27]),
        .b(stage0_col86[28]),
        .c_in(stage0_col86[29]),
        .s(fa_s0_c86_n581_s),
        .c_out(fa_s0_c86_n581_c)
    );

    fa fa_s0_c86_n582 (
        .a(stage0_col86[30]),
        .b(stage0_col86[31]),
        .c_in(stage0_col86[32]),
        .s(fa_s0_c86_n582_s),
        .c_out(fa_s0_c86_n582_c)
    );

    fa fa_s0_c87_n583 (
        .a(stage0_col87[0]),
        .b(stage0_col87[1]),
        .c_in(stage0_col87[2]),
        .s(fa_s0_c87_n583_s),
        .c_out(fa_s0_c87_n583_c)
    );

    fa fa_s0_c87_n584 (
        .a(stage0_col87[3]),
        .b(stage0_col87[4]),
        .c_in(stage0_col87[5]),
        .s(fa_s0_c87_n584_s),
        .c_out(fa_s0_c87_n584_c)
    );

    fa fa_s0_c87_n585 (
        .a(stage0_col87[6]),
        .b(stage0_col87[7]),
        .c_in(stage0_col87[8]),
        .s(fa_s0_c87_n585_s),
        .c_out(fa_s0_c87_n585_c)
    );

    fa fa_s0_c87_n586 (
        .a(stage0_col87[9]),
        .b(stage0_col87[10]),
        .c_in(stage0_col87[11]),
        .s(fa_s0_c87_n586_s),
        .c_out(fa_s0_c87_n586_c)
    );

    fa fa_s0_c87_n587 (
        .a(stage0_col87[12]),
        .b(stage0_col87[13]),
        .c_in(stage0_col87[14]),
        .s(fa_s0_c87_n587_s),
        .c_out(fa_s0_c87_n587_c)
    );

    fa fa_s0_c87_n588 (
        .a(stage0_col87[15]),
        .b(stage0_col87[16]),
        .c_in(stage0_col87[17]),
        .s(fa_s0_c87_n588_s),
        .c_out(fa_s0_c87_n588_c)
    );

    fa fa_s0_c87_n589 (
        .a(stage0_col87[18]),
        .b(stage0_col87[19]),
        .c_in(stage0_col87[20]),
        .s(fa_s0_c87_n589_s),
        .c_out(fa_s0_c87_n589_c)
    );

    fa fa_s0_c87_n590 (
        .a(stage0_col87[21]),
        .b(stage0_col87[22]),
        .c_in(stage0_col87[23]),
        .s(fa_s0_c87_n590_s),
        .c_out(fa_s0_c87_n590_c)
    );

    fa fa_s0_c87_n591 (
        .a(stage0_col87[24]),
        .b(stage0_col87[25]),
        .c_in(stage0_col87[26]),
        .s(fa_s0_c87_n591_s),
        .c_out(fa_s0_c87_n591_c)
    );

    fa fa_s0_c87_n592 (
        .a(stage0_col87[27]),
        .b(stage0_col87[28]),
        .c_in(stage0_col87[29]),
        .s(fa_s0_c87_n592_s),
        .c_out(fa_s0_c87_n592_c)
    );

    fa fa_s0_c88_n593 (
        .a(stage0_col88[0]),
        .b(stage0_col88[1]),
        .c_in(stage0_col88[2]),
        .s(fa_s0_c88_n593_s),
        .c_out(fa_s0_c88_n593_c)
    );

    fa fa_s0_c88_n594 (
        .a(stage0_col88[3]),
        .b(stage0_col88[4]),
        .c_in(stage0_col88[5]),
        .s(fa_s0_c88_n594_s),
        .c_out(fa_s0_c88_n594_c)
    );

    fa fa_s0_c88_n595 (
        .a(stage0_col88[6]),
        .b(stage0_col88[7]),
        .c_in(stage0_col88[8]),
        .s(fa_s0_c88_n595_s),
        .c_out(fa_s0_c88_n595_c)
    );

    fa fa_s0_c88_n596 (
        .a(stage0_col88[9]),
        .b(stage0_col88[10]),
        .c_in(stage0_col88[11]),
        .s(fa_s0_c88_n596_s),
        .c_out(fa_s0_c88_n596_c)
    );

    fa fa_s0_c88_n597 (
        .a(stage0_col88[12]),
        .b(stage0_col88[13]),
        .c_in(stage0_col88[14]),
        .s(fa_s0_c88_n597_s),
        .c_out(fa_s0_c88_n597_c)
    );

    fa fa_s0_c88_n598 (
        .a(stage0_col88[15]),
        .b(stage0_col88[16]),
        .c_in(stage0_col88[17]),
        .s(fa_s0_c88_n598_s),
        .c_out(fa_s0_c88_n598_c)
    );

    fa fa_s0_c88_n599 (
        .a(stage0_col88[18]),
        .b(stage0_col88[19]),
        .c_in(stage0_col88[20]),
        .s(fa_s0_c88_n599_s),
        .c_out(fa_s0_c88_n599_c)
    );

    fa fa_s0_c88_n600 (
        .a(stage0_col88[21]),
        .b(stage0_col88[22]),
        .c_in(stage0_col88[23]),
        .s(fa_s0_c88_n600_s),
        .c_out(fa_s0_c88_n600_c)
    );

    fa fa_s0_c88_n601 (
        .a(stage0_col88[24]),
        .b(stage0_col88[25]),
        .c_in(stage0_col88[26]),
        .s(fa_s0_c88_n601_s),
        .c_out(fa_s0_c88_n601_c)
    );

    fa fa_s0_c88_n602 (
        .a(stage0_col88[27]),
        .b(stage0_col88[28]),
        .c_in(stage0_col88[29]),
        .s(fa_s0_c88_n602_s),
        .c_out(fa_s0_c88_n602_c)
    );

    fa fa_s0_c88_n603 (
        .a(stage0_col88[30]),
        .b(stage0_col88[31]),
        .c_in(stage0_col88[32]),
        .s(fa_s0_c88_n603_s),
        .c_out(fa_s0_c88_n603_c)
    );

    fa fa_s0_c89_n604 (
        .a(stage0_col89[0]),
        .b(stage0_col89[1]),
        .c_in(stage0_col89[2]),
        .s(fa_s0_c89_n604_s),
        .c_out(fa_s0_c89_n604_c)
    );

    fa fa_s0_c89_n605 (
        .a(stage0_col89[3]),
        .b(stage0_col89[4]),
        .c_in(stage0_col89[5]),
        .s(fa_s0_c89_n605_s),
        .c_out(fa_s0_c89_n605_c)
    );

    fa fa_s0_c89_n606 (
        .a(stage0_col89[6]),
        .b(stage0_col89[7]),
        .c_in(stage0_col89[8]),
        .s(fa_s0_c89_n606_s),
        .c_out(fa_s0_c89_n606_c)
    );

    fa fa_s0_c89_n607 (
        .a(stage0_col89[9]),
        .b(stage0_col89[10]),
        .c_in(stage0_col89[11]),
        .s(fa_s0_c89_n607_s),
        .c_out(fa_s0_c89_n607_c)
    );

    fa fa_s0_c89_n608 (
        .a(stage0_col89[12]),
        .b(stage0_col89[13]),
        .c_in(stage0_col89[14]),
        .s(fa_s0_c89_n608_s),
        .c_out(fa_s0_c89_n608_c)
    );

    fa fa_s0_c89_n609 (
        .a(stage0_col89[15]),
        .b(stage0_col89[16]),
        .c_in(stage0_col89[17]),
        .s(fa_s0_c89_n609_s),
        .c_out(fa_s0_c89_n609_c)
    );

    fa fa_s0_c89_n610 (
        .a(stage0_col89[18]),
        .b(stage0_col89[19]),
        .c_in(stage0_col89[20]),
        .s(fa_s0_c89_n610_s),
        .c_out(fa_s0_c89_n610_c)
    );

    fa fa_s0_c89_n611 (
        .a(stage0_col89[21]),
        .b(stage0_col89[22]),
        .c_in(stage0_col89[23]),
        .s(fa_s0_c89_n611_s),
        .c_out(fa_s0_c89_n611_c)
    );

    fa fa_s0_c89_n612 (
        .a(stage0_col89[24]),
        .b(stage0_col89[25]),
        .c_in(stage0_col89[26]),
        .s(fa_s0_c89_n612_s),
        .c_out(fa_s0_c89_n612_c)
    );

    fa fa_s0_c89_n613 (
        .a(stage0_col89[27]),
        .b(stage0_col89[28]),
        .c_in(stage0_col89[29]),
        .s(fa_s0_c89_n613_s),
        .c_out(fa_s0_c89_n613_c)
    );

    fa fa_s0_c90_n614 (
        .a(stage0_col90[0]),
        .b(stage0_col90[1]),
        .c_in(stage0_col90[2]),
        .s(fa_s0_c90_n614_s),
        .c_out(fa_s0_c90_n614_c)
    );

    fa fa_s0_c90_n615 (
        .a(stage0_col90[3]),
        .b(stage0_col90[4]),
        .c_in(stage0_col90[5]),
        .s(fa_s0_c90_n615_s),
        .c_out(fa_s0_c90_n615_c)
    );

    fa fa_s0_c90_n616 (
        .a(stage0_col90[6]),
        .b(stage0_col90[7]),
        .c_in(stage0_col90[8]),
        .s(fa_s0_c90_n616_s),
        .c_out(fa_s0_c90_n616_c)
    );

    fa fa_s0_c90_n617 (
        .a(stage0_col90[9]),
        .b(stage0_col90[10]),
        .c_in(stage0_col90[11]),
        .s(fa_s0_c90_n617_s),
        .c_out(fa_s0_c90_n617_c)
    );

    fa fa_s0_c90_n618 (
        .a(stage0_col90[12]),
        .b(stage0_col90[13]),
        .c_in(stage0_col90[14]),
        .s(fa_s0_c90_n618_s),
        .c_out(fa_s0_c90_n618_c)
    );

    fa fa_s0_c90_n619 (
        .a(stage0_col90[15]),
        .b(stage0_col90[16]),
        .c_in(stage0_col90[17]),
        .s(fa_s0_c90_n619_s),
        .c_out(fa_s0_c90_n619_c)
    );

    fa fa_s0_c90_n620 (
        .a(stage0_col90[18]),
        .b(stage0_col90[19]),
        .c_in(stage0_col90[20]),
        .s(fa_s0_c90_n620_s),
        .c_out(fa_s0_c90_n620_c)
    );

    fa fa_s0_c90_n621 (
        .a(stage0_col90[21]),
        .b(stage0_col90[22]),
        .c_in(stage0_col90[23]),
        .s(fa_s0_c90_n621_s),
        .c_out(fa_s0_c90_n621_c)
    );

    fa fa_s0_c90_n622 (
        .a(stage0_col90[24]),
        .b(stage0_col90[25]),
        .c_in(stage0_col90[26]),
        .s(fa_s0_c90_n622_s),
        .c_out(fa_s0_c90_n622_c)
    );

    fa fa_s0_c90_n623 (
        .a(stage0_col90[27]),
        .b(stage0_col90[28]),
        .c_in(stage0_col90[29]),
        .s(fa_s0_c90_n623_s),
        .c_out(fa_s0_c90_n623_c)
    );

    fa fa_s0_c90_n624 (
        .a(stage0_col90[30]),
        .b(stage0_col90[31]),
        .c_in(stage0_col90[32]),
        .s(fa_s0_c90_n624_s),
        .c_out(fa_s0_c90_n624_c)
    );

    fa fa_s0_c91_n625 (
        .a(stage0_col91[0]),
        .b(stage0_col91[1]),
        .c_in(stage0_col91[2]),
        .s(fa_s0_c91_n625_s),
        .c_out(fa_s0_c91_n625_c)
    );

    fa fa_s0_c91_n626 (
        .a(stage0_col91[3]),
        .b(stage0_col91[4]),
        .c_in(stage0_col91[5]),
        .s(fa_s0_c91_n626_s),
        .c_out(fa_s0_c91_n626_c)
    );

    fa fa_s0_c91_n627 (
        .a(stage0_col91[6]),
        .b(stage0_col91[7]),
        .c_in(stage0_col91[8]),
        .s(fa_s0_c91_n627_s),
        .c_out(fa_s0_c91_n627_c)
    );

    fa fa_s0_c91_n628 (
        .a(stage0_col91[9]),
        .b(stage0_col91[10]),
        .c_in(stage0_col91[11]),
        .s(fa_s0_c91_n628_s),
        .c_out(fa_s0_c91_n628_c)
    );

    fa fa_s0_c91_n629 (
        .a(stage0_col91[12]),
        .b(stage0_col91[13]),
        .c_in(stage0_col91[14]),
        .s(fa_s0_c91_n629_s),
        .c_out(fa_s0_c91_n629_c)
    );

    fa fa_s0_c91_n630 (
        .a(stage0_col91[15]),
        .b(stage0_col91[16]),
        .c_in(stage0_col91[17]),
        .s(fa_s0_c91_n630_s),
        .c_out(fa_s0_c91_n630_c)
    );

    fa fa_s0_c91_n631 (
        .a(stage0_col91[18]),
        .b(stage0_col91[19]),
        .c_in(stage0_col91[20]),
        .s(fa_s0_c91_n631_s),
        .c_out(fa_s0_c91_n631_c)
    );

    fa fa_s0_c91_n632 (
        .a(stage0_col91[21]),
        .b(stage0_col91[22]),
        .c_in(stage0_col91[23]),
        .s(fa_s0_c91_n632_s),
        .c_out(fa_s0_c91_n632_c)
    );

    fa fa_s0_c91_n633 (
        .a(stage0_col91[24]),
        .b(stage0_col91[25]),
        .c_in(stage0_col91[26]),
        .s(fa_s0_c91_n633_s),
        .c_out(fa_s0_c91_n633_c)
    );

    fa fa_s0_c91_n634 (
        .a(stage0_col91[27]),
        .b(stage0_col91[28]),
        .c_in(stage0_col91[29]),
        .s(fa_s0_c91_n634_s),
        .c_out(fa_s0_c91_n634_c)
    );

    fa fa_s0_c92_n635 (
        .a(stage0_col92[0]),
        .b(stage0_col92[1]),
        .c_in(stage0_col92[2]),
        .s(fa_s0_c92_n635_s),
        .c_out(fa_s0_c92_n635_c)
    );

    fa fa_s0_c92_n636 (
        .a(stage0_col92[3]),
        .b(stage0_col92[4]),
        .c_in(stage0_col92[5]),
        .s(fa_s0_c92_n636_s),
        .c_out(fa_s0_c92_n636_c)
    );

    fa fa_s0_c92_n637 (
        .a(stage0_col92[6]),
        .b(stage0_col92[7]),
        .c_in(stage0_col92[8]),
        .s(fa_s0_c92_n637_s),
        .c_out(fa_s0_c92_n637_c)
    );

    fa fa_s0_c92_n638 (
        .a(stage0_col92[9]),
        .b(stage0_col92[10]),
        .c_in(stage0_col92[11]),
        .s(fa_s0_c92_n638_s),
        .c_out(fa_s0_c92_n638_c)
    );

    fa fa_s0_c92_n639 (
        .a(stage0_col92[12]),
        .b(stage0_col92[13]),
        .c_in(stage0_col92[14]),
        .s(fa_s0_c92_n639_s),
        .c_out(fa_s0_c92_n639_c)
    );

    fa fa_s0_c92_n640 (
        .a(stage0_col92[15]),
        .b(stage0_col92[16]),
        .c_in(stage0_col92[17]),
        .s(fa_s0_c92_n640_s),
        .c_out(fa_s0_c92_n640_c)
    );

    fa fa_s0_c92_n641 (
        .a(stage0_col92[18]),
        .b(stage0_col92[19]),
        .c_in(stage0_col92[20]),
        .s(fa_s0_c92_n641_s),
        .c_out(fa_s0_c92_n641_c)
    );

    fa fa_s0_c92_n642 (
        .a(stage0_col92[21]),
        .b(stage0_col92[22]),
        .c_in(stage0_col92[23]),
        .s(fa_s0_c92_n642_s),
        .c_out(fa_s0_c92_n642_c)
    );

    fa fa_s0_c92_n643 (
        .a(stage0_col92[24]),
        .b(stage0_col92[25]),
        .c_in(stage0_col92[26]),
        .s(fa_s0_c92_n643_s),
        .c_out(fa_s0_c92_n643_c)
    );

    fa fa_s0_c92_n644 (
        .a(stage0_col92[27]),
        .b(stage0_col92[28]),
        .c_in(stage0_col92[29]),
        .s(fa_s0_c92_n644_s),
        .c_out(fa_s0_c92_n644_c)
    );

    fa fa_s0_c92_n645 (
        .a(stage0_col92[30]),
        .b(stage0_col92[31]),
        .c_in(stage0_col92[32]),
        .s(fa_s0_c92_n645_s),
        .c_out(fa_s0_c92_n645_c)
    );

    fa fa_s0_c93_n646 (
        .a(stage0_col93[0]),
        .b(stage0_col93[1]),
        .c_in(stage0_col93[2]),
        .s(fa_s0_c93_n646_s),
        .c_out(fa_s0_c93_n646_c)
    );

    fa fa_s0_c93_n647 (
        .a(stage0_col93[3]),
        .b(stage0_col93[4]),
        .c_in(stage0_col93[5]),
        .s(fa_s0_c93_n647_s),
        .c_out(fa_s0_c93_n647_c)
    );

    fa fa_s0_c93_n648 (
        .a(stage0_col93[6]),
        .b(stage0_col93[7]),
        .c_in(stage0_col93[8]),
        .s(fa_s0_c93_n648_s),
        .c_out(fa_s0_c93_n648_c)
    );

    fa fa_s0_c93_n649 (
        .a(stage0_col93[9]),
        .b(stage0_col93[10]),
        .c_in(stage0_col93[11]),
        .s(fa_s0_c93_n649_s),
        .c_out(fa_s0_c93_n649_c)
    );

    fa fa_s0_c93_n650 (
        .a(stage0_col93[12]),
        .b(stage0_col93[13]),
        .c_in(stage0_col93[14]),
        .s(fa_s0_c93_n650_s),
        .c_out(fa_s0_c93_n650_c)
    );

    fa fa_s0_c93_n651 (
        .a(stage0_col93[15]),
        .b(stage0_col93[16]),
        .c_in(stage0_col93[17]),
        .s(fa_s0_c93_n651_s),
        .c_out(fa_s0_c93_n651_c)
    );

    fa fa_s0_c93_n652 (
        .a(stage0_col93[18]),
        .b(stage0_col93[19]),
        .c_in(stage0_col93[20]),
        .s(fa_s0_c93_n652_s),
        .c_out(fa_s0_c93_n652_c)
    );

    fa fa_s0_c93_n653 (
        .a(stage0_col93[21]),
        .b(stage0_col93[22]),
        .c_in(stage0_col93[23]),
        .s(fa_s0_c93_n653_s),
        .c_out(fa_s0_c93_n653_c)
    );

    fa fa_s0_c93_n654 (
        .a(stage0_col93[24]),
        .b(stage0_col93[25]),
        .c_in(stage0_col93[26]),
        .s(fa_s0_c93_n654_s),
        .c_out(fa_s0_c93_n654_c)
    );

    fa fa_s0_c93_n655 (
        .a(stage0_col93[27]),
        .b(stage0_col93[28]),
        .c_in(stage0_col93[29]),
        .s(fa_s0_c93_n655_s),
        .c_out(fa_s0_c93_n655_c)
    );

    fa fa_s0_c94_n656 (
        .a(stage0_col94[0]),
        .b(stage0_col94[1]),
        .c_in(stage0_col94[2]),
        .s(fa_s0_c94_n656_s),
        .c_out(fa_s0_c94_n656_c)
    );

    fa fa_s0_c94_n657 (
        .a(stage0_col94[3]),
        .b(stage0_col94[4]),
        .c_in(stage0_col94[5]),
        .s(fa_s0_c94_n657_s),
        .c_out(fa_s0_c94_n657_c)
    );

    fa fa_s0_c94_n658 (
        .a(stage0_col94[6]),
        .b(stage0_col94[7]),
        .c_in(stage0_col94[8]),
        .s(fa_s0_c94_n658_s),
        .c_out(fa_s0_c94_n658_c)
    );

    fa fa_s0_c94_n659 (
        .a(stage0_col94[9]),
        .b(stage0_col94[10]),
        .c_in(stage0_col94[11]),
        .s(fa_s0_c94_n659_s),
        .c_out(fa_s0_c94_n659_c)
    );

    fa fa_s0_c94_n660 (
        .a(stage0_col94[12]),
        .b(stage0_col94[13]),
        .c_in(stage0_col94[14]),
        .s(fa_s0_c94_n660_s),
        .c_out(fa_s0_c94_n660_c)
    );

    fa fa_s0_c94_n661 (
        .a(stage0_col94[15]),
        .b(stage0_col94[16]),
        .c_in(stage0_col94[17]),
        .s(fa_s0_c94_n661_s),
        .c_out(fa_s0_c94_n661_c)
    );

    fa fa_s0_c94_n662 (
        .a(stage0_col94[18]),
        .b(stage0_col94[19]),
        .c_in(stage0_col94[20]),
        .s(fa_s0_c94_n662_s),
        .c_out(fa_s0_c94_n662_c)
    );

    fa fa_s0_c94_n663 (
        .a(stage0_col94[21]),
        .b(stage0_col94[22]),
        .c_in(stage0_col94[23]),
        .s(fa_s0_c94_n663_s),
        .c_out(fa_s0_c94_n663_c)
    );

    fa fa_s0_c94_n664 (
        .a(stage0_col94[24]),
        .b(stage0_col94[25]),
        .c_in(stage0_col94[26]),
        .s(fa_s0_c94_n664_s),
        .c_out(fa_s0_c94_n664_c)
    );

    fa fa_s0_c94_n665 (
        .a(stage0_col94[27]),
        .b(stage0_col94[28]),
        .c_in(stage0_col94[29]),
        .s(fa_s0_c94_n665_s),
        .c_out(fa_s0_c94_n665_c)
    );

    fa fa_s0_c94_n666 (
        .a(stage0_col94[30]),
        .b(stage0_col94[31]),
        .c_in(stage0_col94[32]),
        .s(fa_s0_c94_n666_s),
        .c_out(fa_s0_c94_n666_c)
    );

    fa fa_s0_c95_n667 (
        .a(stage0_col95[0]),
        .b(stage0_col95[1]),
        .c_in(stage0_col95[2]),
        .s(fa_s0_c95_n667_s),
        .c_out(fa_s0_c95_n667_c)
    );

    fa fa_s0_c95_n668 (
        .a(stage0_col95[3]),
        .b(stage0_col95[4]),
        .c_in(stage0_col95[5]),
        .s(fa_s0_c95_n668_s),
        .c_out(fa_s0_c95_n668_c)
    );

    fa fa_s0_c95_n669 (
        .a(stage0_col95[6]),
        .b(stage0_col95[7]),
        .c_in(stage0_col95[8]),
        .s(fa_s0_c95_n669_s),
        .c_out(fa_s0_c95_n669_c)
    );

    fa fa_s0_c95_n670 (
        .a(stage0_col95[9]),
        .b(stage0_col95[10]),
        .c_in(stage0_col95[11]),
        .s(fa_s0_c95_n670_s),
        .c_out(fa_s0_c95_n670_c)
    );

    fa fa_s0_c95_n671 (
        .a(stage0_col95[12]),
        .b(stage0_col95[13]),
        .c_in(stage0_col95[14]),
        .s(fa_s0_c95_n671_s),
        .c_out(fa_s0_c95_n671_c)
    );

    fa fa_s0_c95_n672 (
        .a(stage0_col95[15]),
        .b(stage0_col95[16]),
        .c_in(stage0_col95[17]),
        .s(fa_s0_c95_n672_s),
        .c_out(fa_s0_c95_n672_c)
    );

    fa fa_s0_c95_n673 (
        .a(stage0_col95[18]),
        .b(stage0_col95[19]),
        .c_in(stage0_col95[20]),
        .s(fa_s0_c95_n673_s),
        .c_out(fa_s0_c95_n673_c)
    );

    fa fa_s0_c95_n674 (
        .a(stage0_col95[21]),
        .b(stage0_col95[22]),
        .c_in(stage0_col95[23]),
        .s(fa_s0_c95_n674_s),
        .c_out(fa_s0_c95_n674_c)
    );

    fa fa_s0_c95_n675 (
        .a(stage0_col95[24]),
        .b(stage0_col95[25]),
        .c_in(stage0_col95[26]),
        .s(fa_s0_c95_n675_s),
        .c_out(fa_s0_c95_n675_c)
    );

    fa fa_s0_c95_n676 (
        .a(stage0_col95[27]),
        .b(stage0_col95[28]),
        .c_in(stage0_col95[29]),
        .s(fa_s0_c95_n676_s),
        .c_out(fa_s0_c95_n676_c)
    );

    fa fa_s0_c96_n677 (
        .a(stage0_col96[0]),
        .b(stage0_col96[1]),
        .c_in(stage0_col96[2]),
        .s(fa_s0_c96_n677_s),
        .c_out(fa_s0_c96_n677_c)
    );

    fa fa_s0_c96_n678 (
        .a(stage0_col96[3]),
        .b(stage0_col96[4]),
        .c_in(stage0_col96[5]),
        .s(fa_s0_c96_n678_s),
        .c_out(fa_s0_c96_n678_c)
    );

    fa fa_s0_c96_n679 (
        .a(stage0_col96[6]),
        .b(stage0_col96[7]),
        .c_in(stage0_col96[8]),
        .s(fa_s0_c96_n679_s),
        .c_out(fa_s0_c96_n679_c)
    );

    fa fa_s0_c96_n680 (
        .a(stage0_col96[9]),
        .b(stage0_col96[10]),
        .c_in(stage0_col96[11]),
        .s(fa_s0_c96_n680_s),
        .c_out(fa_s0_c96_n680_c)
    );

    fa fa_s0_c96_n681 (
        .a(stage0_col96[12]),
        .b(stage0_col96[13]),
        .c_in(stage0_col96[14]),
        .s(fa_s0_c96_n681_s),
        .c_out(fa_s0_c96_n681_c)
    );

    fa fa_s0_c96_n682 (
        .a(stage0_col96[15]),
        .b(stage0_col96[16]),
        .c_in(stage0_col96[17]),
        .s(fa_s0_c96_n682_s),
        .c_out(fa_s0_c96_n682_c)
    );

    fa fa_s0_c96_n683 (
        .a(stage0_col96[18]),
        .b(stage0_col96[19]),
        .c_in(stage0_col96[20]),
        .s(fa_s0_c96_n683_s),
        .c_out(fa_s0_c96_n683_c)
    );

    fa fa_s0_c96_n684 (
        .a(stage0_col96[21]),
        .b(stage0_col96[22]),
        .c_in(stage0_col96[23]),
        .s(fa_s0_c96_n684_s),
        .c_out(fa_s0_c96_n684_c)
    );

    fa fa_s0_c96_n685 (
        .a(stage0_col96[24]),
        .b(stage0_col96[25]),
        .c_in(stage0_col96[26]),
        .s(fa_s0_c96_n685_s),
        .c_out(fa_s0_c96_n685_c)
    );

    fa fa_s0_c96_n686 (
        .a(stage0_col96[27]),
        .b(stage0_col96[28]),
        .c_in(stage0_col96[29]),
        .s(fa_s0_c96_n686_s),
        .c_out(fa_s0_c96_n686_c)
    );

    fa fa_s0_c96_n687 (
        .a(stage0_col96[30]),
        .b(stage0_col96[31]),
        .c_in(stage0_col96[32]),
        .s(fa_s0_c96_n687_s),
        .c_out(fa_s0_c96_n687_c)
    );

    fa fa_s0_c97_n688 (
        .a(stage0_col97[0]),
        .b(stage0_col97[1]),
        .c_in(stage0_col97[2]),
        .s(fa_s0_c97_n688_s),
        .c_out(fa_s0_c97_n688_c)
    );

    fa fa_s0_c97_n689 (
        .a(stage0_col97[3]),
        .b(stage0_col97[4]),
        .c_in(stage0_col97[5]),
        .s(fa_s0_c97_n689_s),
        .c_out(fa_s0_c97_n689_c)
    );

    fa fa_s0_c97_n690 (
        .a(stage0_col97[6]),
        .b(stage0_col97[7]),
        .c_in(stage0_col97[8]),
        .s(fa_s0_c97_n690_s),
        .c_out(fa_s0_c97_n690_c)
    );

    fa fa_s0_c97_n691 (
        .a(stage0_col97[9]),
        .b(stage0_col97[10]),
        .c_in(stage0_col97[11]),
        .s(fa_s0_c97_n691_s),
        .c_out(fa_s0_c97_n691_c)
    );

    fa fa_s0_c97_n692 (
        .a(stage0_col97[12]),
        .b(stage0_col97[13]),
        .c_in(stage0_col97[14]),
        .s(fa_s0_c97_n692_s),
        .c_out(fa_s0_c97_n692_c)
    );

    fa fa_s0_c97_n693 (
        .a(stage0_col97[15]),
        .b(stage0_col97[16]),
        .c_in(stage0_col97[17]),
        .s(fa_s0_c97_n693_s),
        .c_out(fa_s0_c97_n693_c)
    );

    fa fa_s0_c97_n694 (
        .a(stage0_col97[18]),
        .b(stage0_col97[19]),
        .c_in(stage0_col97[20]),
        .s(fa_s0_c97_n694_s),
        .c_out(fa_s0_c97_n694_c)
    );

    fa fa_s0_c97_n695 (
        .a(stage0_col97[21]),
        .b(stage0_col97[22]),
        .c_in(stage0_col97[23]),
        .s(fa_s0_c97_n695_s),
        .c_out(fa_s0_c97_n695_c)
    );

    fa fa_s0_c97_n696 (
        .a(stage0_col97[24]),
        .b(stage0_col97[25]),
        .c_in(stage0_col97[26]),
        .s(fa_s0_c97_n696_s),
        .c_out(fa_s0_c97_n696_c)
    );

    fa fa_s0_c97_n697 (
        .a(stage0_col97[27]),
        .b(stage0_col97[28]),
        .c_in(stage0_col97[29]),
        .s(fa_s0_c97_n697_s),
        .c_out(fa_s0_c97_n697_c)
    );

    fa fa_s0_c98_n698 (
        .a(stage0_col98[0]),
        .b(stage0_col98[1]),
        .c_in(stage0_col98[2]),
        .s(fa_s0_c98_n698_s),
        .c_out(fa_s0_c98_n698_c)
    );

    fa fa_s0_c98_n699 (
        .a(stage0_col98[3]),
        .b(stage0_col98[4]),
        .c_in(stage0_col98[5]),
        .s(fa_s0_c98_n699_s),
        .c_out(fa_s0_c98_n699_c)
    );

    fa fa_s0_c98_n700 (
        .a(stage0_col98[6]),
        .b(stage0_col98[7]),
        .c_in(stage0_col98[8]),
        .s(fa_s0_c98_n700_s),
        .c_out(fa_s0_c98_n700_c)
    );

    fa fa_s0_c98_n701 (
        .a(stage0_col98[9]),
        .b(stage0_col98[10]),
        .c_in(stage0_col98[11]),
        .s(fa_s0_c98_n701_s),
        .c_out(fa_s0_c98_n701_c)
    );

    fa fa_s0_c98_n702 (
        .a(stage0_col98[12]),
        .b(stage0_col98[13]),
        .c_in(stage0_col98[14]),
        .s(fa_s0_c98_n702_s),
        .c_out(fa_s0_c98_n702_c)
    );

    fa fa_s0_c98_n703 (
        .a(stage0_col98[15]),
        .b(stage0_col98[16]),
        .c_in(stage0_col98[17]),
        .s(fa_s0_c98_n703_s),
        .c_out(fa_s0_c98_n703_c)
    );

    fa fa_s0_c98_n704 (
        .a(stage0_col98[18]),
        .b(stage0_col98[19]),
        .c_in(stage0_col98[20]),
        .s(fa_s0_c98_n704_s),
        .c_out(fa_s0_c98_n704_c)
    );

    fa fa_s0_c98_n705 (
        .a(stage0_col98[21]),
        .b(stage0_col98[22]),
        .c_in(stage0_col98[23]),
        .s(fa_s0_c98_n705_s),
        .c_out(fa_s0_c98_n705_c)
    );

    fa fa_s0_c98_n706 (
        .a(stage0_col98[24]),
        .b(stage0_col98[25]),
        .c_in(stage0_col98[26]),
        .s(fa_s0_c98_n706_s),
        .c_out(fa_s0_c98_n706_c)
    );

    fa fa_s0_c98_n707 (
        .a(stage0_col98[27]),
        .b(stage0_col98[28]),
        .c_in(stage0_col98[29]),
        .s(fa_s0_c98_n707_s),
        .c_out(fa_s0_c98_n707_c)
    );

    fa fa_s0_c98_n708 (
        .a(stage0_col98[30]),
        .b(stage0_col98[31]),
        .c_in(stage0_col98[32]),
        .s(fa_s0_c98_n708_s),
        .c_out(fa_s0_c98_n708_c)
    );

    fa fa_s0_c99_n709 (
        .a(stage0_col99[0]),
        .b(stage0_col99[1]),
        .c_in(stage0_col99[2]),
        .s(fa_s0_c99_n709_s),
        .c_out(fa_s0_c99_n709_c)
    );

    fa fa_s0_c99_n710 (
        .a(stage0_col99[3]),
        .b(stage0_col99[4]),
        .c_in(stage0_col99[5]),
        .s(fa_s0_c99_n710_s),
        .c_out(fa_s0_c99_n710_c)
    );

    fa fa_s0_c99_n711 (
        .a(stage0_col99[6]),
        .b(stage0_col99[7]),
        .c_in(stage0_col99[8]),
        .s(fa_s0_c99_n711_s),
        .c_out(fa_s0_c99_n711_c)
    );

    fa fa_s0_c99_n712 (
        .a(stage0_col99[9]),
        .b(stage0_col99[10]),
        .c_in(stage0_col99[11]),
        .s(fa_s0_c99_n712_s),
        .c_out(fa_s0_c99_n712_c)
    );

    fa fa_s0_c99_n713 (
        .a(stage0_col99[12]),
        .b(stage0_col99[13]),
        .c_in(stage0_col99[14]),
        .s(fa_s0_c99_n713_s),
        .c_out(fa_s0_c99_n713_c)
    );

    fa fa_s0_c99_n714 (
        .a(stage0_col99[15]),
        .b(stage0_col99[16]),
        .c_in(stage0_col99[17]),
        .s(fa_s0_c99_n714_s),
        .c_out(fa_s0_c99_n714_c)
    );

    fa fa_s0_c99_n715 (
        .a(stage0_col99[18]),
        .b(stage0_col99[19]),
        .c_in(stage0_col99[20]),
        .s(fa_s0_c99_n715_s),
        .c_out(fa_s0_c99_n715_c)
    );

    fa fa_s0_c99_n716 (
        .a(stage0_col99[21]),
        .b(stage0_col99[22]),
        .c_in(stage0_col99[23]),
        .s(fa_s0_c99_n716_s),
        .c_out(fa_s0_c99_n716_c)
    );

    fa fa_s0_c99_n717 (
        .a(stage0_col99[24]),
        .b(stage0_col99[25]),
        .c_in(stage0_col99[26]),
        .s(fa_s0_c99_n717_s),
        .c_out(fa_s0_c99_n717_c)
    );

    fa fa_s0_c99_n718 (
        .a(stage0_col99[27]),
        .b(stage0_col99[28]),
        .c_in(stage0_col99[29]),
        .s(fa_s0_c99_n718_s),
        .c_out(fa_s0_c99_n718_c)
    );

    fa fa_s0_c100_n719 (
        .a(stage0_col100[0]),
        .b(stage0_col100[1]),
        .c_in(stage0_col100[2]),
        .s(fa_s0_c100_n719_s),
        .c_out(fa_s0_c100_n719_c)
    );

    fa fa_s0_c100_n720 (
        .a(stage0_col100[3]),
        .b(stage0_col100[4]),
        .c_in(stage0_col100[5]),
        .s(fa_s0_c100_n720_s),
        .c_out(fa_s0_c100_n720_c)
    );

    fa fa_s0_c100_n721 (
        .a(stage0_col100[6]),
        .b(stage0_col100[7]),
        .c_in(stage0_col100[8]),
        .s(fa_s0_c100_n721_s),
        .c_out(fa_s0_c100_n721_c)
    );

    fa fa_s0_c100_n722 (
        .a(stage0_col100[9]),
        .b(stage0_col100[10]),
        .c_in(stage0_col100[11]),
        .s(fa_s0_c100_n722_s),
        .c_out(fa_s0_c100_n722_c)
    );

    fa fa_s0_c100_n723 (
        .a(stage0_col100[12]),
        .b(stage0_col100[13]),
        .c_in(stage0_col100[14]),
        .s(fa_s0_c100_n723_s),
        .c_out(fa_s0_c100_n723_c)
    );

    fa fa_s0_c100_n724 (
        .a(stage0_col100[15]),
        .b(stage0_col100[16]),
        .c_in(stage0_col100[17]),
        .s(fa_s0_c100_n724_s),
        .c_out(fa_s0_c100_n724_c)
    );

    fa fa_s0_c100_n725 (
        .a(stage0_col100[18]),
        .b(stage0_col100[19]),
        .c_in(stage0_col100[20]),
        .s(fa_s0_c100_n725_s),
        .c_out(fa_s0_c100_n725_c)
    );

    fa fa_s0_c100_n726 (
        .a(stage0_col100[21]),
        .b(stage0_col100[22]),
        .c_in(stage0_col100[23]),
        .s(fa_s0_c100_n726_s),
        .c_out(fa_s0_c100_n726_c)
    );

    fa fa_s0_c100_n727 (
        .a(stage0_col100[24]),
        .b(stage0_col100[25]),
        .c_in(stage0_col100[26]),
        .s(fa_s0_c100_n727_s),
        .c_out(fa_s0_c100_n727_c)
    );

    fa fa_s0_c100_n728 (
        .a(stage0_col100[27]),
        .b(stage0_col100[28]),
        .c_in(stage0_col100[29]),
        .s(fa_s0_c100_n728_s),
        .c_out(fa_s0_c100_n728_c)
    );

    fa fa_s0_c100_n729 (
        .a(stage0_col100[30]),
        .b(stage0_col100[31]),
        .c_in(stage0_col100[32]),
        .s(fa_s0_c100_n729_s),
        .c_out(fa_s0_c100_n729_c)
    );

    fa fa_s0_c101_n730 (
        .a(stage0_col101[0]),
        .b(stage0_col101[1]),
        .c_in(stage0_col101[2]),
        .s(fa_s0_c101_n730_s),
        .c_out(fa_s0_c101_n730_c)
    );

    fa fa_s0_c101_n731 (
        .a(stage0_col101[3]),
        .b(stage0_col101[4]),
        .c_in(stage0_col101[5]),
        .s(fa_s0_c101_n731_s),
        .c_out(fa_s0_c101_n731_c)
    );

    fa fa_s0_c101_n732 (
        .a(stage0_col101[6]),
        .b(stage0_col101[7]),
        .c_in(stage0_col101[8]),
        .s(fa_s0_c101_n732_s),
        .c_out(fa_s0_c101_n732_c)
    );

    fa fa_s0_c101_n733 (
        .a(stage0_col101[9]),
        .b(stage0_col101[10]),
        .c_in(stage0_col101[11]),
        .s(fa_s0_c101_n733_s),
        .c_out(fa_s0_c101_n733_c)
    );

    fa fa_s0_c101_n734 (
        .a(stage0_col101[12]),
        .b(stage0_col101[13]),
        .c_in(stage0_col101[14]),
        .s(fa_s0_c101_n734_s),
        .c_out(fa_s0_c101_n734_c)
    );

    fa fa_s0_c101_n735 (
        .a(stage0_col101[15]),
        .b(stage0_col101[16]),
        .c_in(stage0_col101[17]),
        .s(fa_s0_c101_n735_s),
        .c_out(fa_s0_c101_n735_c)
    );

    fa fa_s0_c101_n736 (
        .a(stage0_col101[18]),
        .b(stage0_col101[19]),
        .c_in(stage0_col101[20]),
        .s(fa_s0_c101_n736_s),
        .c_out(fa_s0_c101_n736_c)
    );

    fa fa_s0_c101_n737 (
        .a(stage0_col101[21]),
        .b(stage0_col101[22]),
        .c_in(stage0_col101[23]),
        .s(fa_s0_c101_n737_s),
        .c_out(fa_s0_c101_n737_c)
    );

    fa fa_s0_c101_n738 (
        .a(stage0_col101[24]),
        .b(stage0_col101[25]),
        .c_in(stage0_col101[26]),
        .s(fa_s0_c101_n738_s),
        .c_out(fa_s0_c101_n738_c)
    );

    fa fa_s0_c101_n739 (
        .a(stage0_col101[27]),
        .b(stage0_col101[28]),
        .c_in(stage0_col101[29]),
        .s(fa_s0_c101_n739_s),
        .c_out(fa_s0_c101_n739_c)
    );

    fa fa_s0_c102_n740 (
        .a(stage0_col102[0]),
        .b(stage0_col102[1]),
        .c_in(stage0_col102[2]),
        .s(fa_s0_c102_n740_s),
        .c_out(fa_s0_c102_n740_c)
    );

    fa fa_s0_c102_n741 (
        .a(stage0_col102[3]),
        .b(stage0_col102[4]),
        .c_in(stage0_col102[5]),
        .s(fa_s0_c102_n741_s),
        .c_out(fa_s0_c102_n741_c)
    );

    fa fa_s0_c102_n742 (
        .a(stage0_col102[6]),
        .b(stage0_col102[7]),
        .c_in(stage0_col102[8]),
        .s(fa_s0_c102_n742_s),
        .c_out(fa_s0_c102_n742_c)
    );

    fa fa_s0_c102_n743 (
        .a(stage0_col102[9]),
        .b(stage0_col102[10]),
        .c_in(stage0_col102[11]),
        .s(fa_s0_c102_n743_s),
        .c_out(fa_s0_c102_n743_c)
    );

    fa fa_s0_c102_n744 (
        .a(stage0_col102[12]),
        .b(stage0_col102[13]),
        .c_in(stage0_col102[14]),
        .s(fa_s0_c102_n744_s),
        .c_out(fa_s0_c102_n744_c)
    );

    fa fa_s0_c102_n745 (
        .a(stage0_col102[15]),
        .b(stage0_col102[16]),
        .c_in(stage0_col102[17]),
        .s(fa_s0_c102_n745_s),
        .c_out(fa_s0_c102_n745_c)
    );

    fa fa_s0_c102_n746 (
        .a(stage0_col102[18]),
        .b(stage0_col102[19]),
        .c_in(stage0_col102[20]),
        .s(fa_s0_c102_n746_s),
        .c_out(fa_s0_c102_n746_c)
    );

    fa fa_s0_c102_n747 (
        .a(stage0_col102[21]),
        .b(stage0_col102[22]),
        .c_in(stage0_col102[23]),
        .s(fa_s0_c102_n747_s),
        .c_out(fa_s0_c102_n747_c)
    );

    fa fa_s0_c102_n748 (
        .a(stage0_col102[24]),
        .b(stage0_col102[25]),
        .c_in(stage0_col102[26]),
        .s(fa_s0_c102_n748_s),
        .c_out(fa_s0_c102_n748_c)
    );

    fa fa_s0_c102_n749 (
        .a(stage0_col102[27]),
        .b(stage0_col102[28]),
        .c_in(stage0_col102[29]),
        .s(fa_s0_c102_n749_s),
        .c_out(fa_s0_c102_n749_c)
    );

    fa fa_s0_c102_n750 (
        .a(stage0_col102[30]),
        .b(stage0_col102[31]),
        .c_in(stage0_col102[32]),
        .s(fa_s0_c102_n750_s),
        .c_out(fa_s0_c102_n750_c)
    );

    fa fa_s0_c103_n751 (
        .a(stage0_col103[0]),
        .b(stage0_col103[1]),
        .c_in(stage0_col103[2]),
        .s(fa_s0_c103_n751_s),
        .c_out(fa_s0_c103_n751_c)
    );

    fa fa_s0_c103_n752 (
        .a(stage0_col103[3]),
        .b(stage0_col103[4]),
        .c_in(stage0_col103[5]),
        .s(fa_s0_c103_n752_s),
        .c_out(fa_s0_c103_n752_c)
    );

    fa fa_s0_c103_n753 (
        .a(stage0_col103[6]),
        .b(stage0_col103[7]),
        .c_in(stage0_col103[8]),
        .s(fa_s0_c103_n753_s),
        .c_out(fa_s0_c103_n753_c)
    );

    fa fa_s0_c103_n754 (
        .a(stage0_col103[9]),
        .b(stage0_col103[10]),
        .c_in(stage0_col103[11]),
        .s(fa_s0_c103_n754_s),
        .c_out(fa_s0_c103_n754_c)
    );

    fa fa_s0_c103_n755 (
        .a(stage0_col103[12]),
        .b(stage0_col103[13]),
        .c_in(stage0_col103[14]),
        .s(fa_s0_c103_n755_s),
        .c_out(fa_s0_c103_n755_c)
    );

    fa fa_s0_c103_n756 (
        .a(stage0_col103[15]),
        .b(stage0_col103[16]),
        .c_in(stage0_col103[17]),
        .s(fa_s0_c103_n756_s),
        .c_out(fa_s0_c103_n756_c)
    );

    fa fa_s0_c103_n757 (
        .a(stage0_col103[18]),
        .b(stage0_col103[19]),
        .c_in(stage0_col103[20]),
        .s(fa_s0_c103_n757_s),
        .c_out(fa_s0_c103_n757_c)
    );

    fa fa_s0_c103_n758 (
        .a(stage0_col103[21]),
        .b(stage0_col103[22]),
        .c_in(stage0_col103[23]),
        .s(fa_s0_c103_n758_s),
        .c_out(fa_s0_c103_n758_c)
    );

    fa fa_s0_c103_n759 (
        .a(stage0_col103[24]),
        .b(stage0_col103[25]),
        .c_in(stage0_col103[26]),
        .s(fa_s0_c103_n759_s),
        .c_out(fa_s0_c103_n759_c)
    );

    fa fa_s0_c103_n760 (
        .a(stage0_col103[27]),
        .b(stage0_col103[28]),
        .c_in(stage0_col103[29]),
        .s(fa_s0_c103_n760_s),
        .c_out(fa_s0_c103_n760_c)
    );

    fa fa_s0_c104_n761 (
        .a(stage0_col104[0]),
        .b(stage0_col104[1]),
        .c_in(stage0_col104[2]),
        .s(fa_s0_c104_n761_s),
        .c_out(fa_s0_c104_n761_c)
    );

    fa fa_s0_c104_n762 (
        .a(stage0_col104[3]),
        .b(stage0_col104[4]),
        .c_in(stage0_col104[5]),
        .s(fa_s0_c104_n762_s),
        .c_out(fa_s0_c104_n762_c)
    );

    fa fa_s0_c104_n763 (
        .a(stage0_col104[6]),
        .b(stage0_col104[7]),
        .c_in(stage0_col104[8]),
        .s(fa_s0_c104_n763_s),
        .c_out(fa_s0_c104_n763_c)
    );

    fa fa_s0_c104_n764 (
        .a(stage0_col104[9]),
        .b(stage0_col104[10]),
        .c_in(stage0_col104[11]),
        .s(fa_s0_c104_n764_s),
        .c_out(fa_s0_c104_n764_c)
    );

    fa fa_s0_c104_n765 (
        .a(stage0_col104[12]),
        .b(stage0_col104[13]),
        .c_in(stage0_col104[14]),
        .s(fa_s0_c104_n765_s),
        .c_out(fa_s0_c104_n765_c)
    );

    fa fa_s0_c104_n766 (
        .a(stage0_col104[15]),
        .b(stage0_col104[16]),
        .c_in(stage0_col104[17]),
        .s(fa_s0_c104_n766_s),
        .c_out(fa_s0_c104_n766_c)
    );

    fa fa_s0_c104_n767 (
        .a(stage0_col104[18]),
        .b(stage0_col104[19]),
        .c_in(stage0_col104[20]),
        .s(fa_s0_c104_n767_s),
        .c_out(fa_s0_c104_n767_c)
    );

    fa fa_s0_c104_n768 (
        .a(stage0_col104[21]),
        .b(stage0_col104[22]),
        .c_in(stage0_col104[23]),
        .s(fa_s0_c104_n768_s),
        .c_out(fa_s0_c104_n768_c)
    );

    fa fa_s0_c104_n769 (
        .a(stage0_col104[24]),
        .b(stage0_col104[25]),
        .c_in(stage0_col104[26]),
        .s(fa_s0_c104_n769_s),
        .c_out(fa_s0_c104_n769_c)
    );

    fa fa_s0_c104_n770 (
        .a(stage0_col104[27]),
        .b(stage0_col104[28]),
        .c_in(stage0_col104[29]),
        .s(fa_s0_c104_n770_s),
        .c_out(fa_s0_c104_n770_c)
    );

    fa fa_s0_c104_n771 (
        .a(stage0_col104[30]),
        .b(stage0_col104[31]),
        .c_in(stage0_col104[32]),
        .s(fa_s0_c104_n771_s),
        .c_out(fa_s0_c104_n771_c)
    );

    fa fa_s0_c105_n772 (
        .a(stage0_col105[0]),
        .b(stage0_col105[1]),
        .c_in(stage0_col105[2]),
        .s(fa_s0_c105_n772_s),
        .c_out(fa_s0_c105_n772_c)
    );

    fa fa_s0_c105_n773 (
        .a(stage0_col105[3]),
        .b(stage0_col105[4]),
        .c_in(stage0_col105[5]),
        .s(fa_s0_c105_n773_s),
        .c_out(fa_s0_c105_n773_c)
    );

    fa fa_s0_c105_n774 (
        .a(stage0_col105[6]),
        .b(stage0_col105[7]),
        .c_in(stage0_col105[8]),
        .s(fa_s0_c105_n774_s),
        .c_out(fa_s0_c105_n774_c)
    );

    fa fa_s0_c105_n775 (
        .a(stage0_col105[9]),
        .b(stage0_col105[10]),
        .c_in(stage0_col105[11]),
        .s(fa_s0_c105_n775_s),
        .c_out(fa_s0_c105_n775_c)
    );

    fa fa_s0_c105_n776 (
        .a(stage0_col105[12]),
        .b(stage0_col105[13]),
        .c_in(stage0_col105[14]),
        .s(fa_s0_c105_n776_s),
        .c_out(fa_s0_c105_n776_c)
    );

    fa fa_s0_c105_n777 (
        .a(stage0_col105[15]),
        .b(stage0_col105[16]),
        .c_in(stage0_col105[17]),
        .s(fa_s0_c105_n777_s),
        .c_out(fa_s0_c105_n777_c)
    );

    fa fa_s0_c105_n778 (
        .a(stage0_col105[18]),
        .b(stage0_col105[19]),
        .c_in(stage0_col105[20]),
        .s(fa_s0_c105_n778_s),
        .c_out(fa_s0_c105_n778_c)
    );

    fa fa_s0_c105_n779 (
        .a(stage0_col105[21]),
        .b(stage0_col105[22]),
        .c_in(stage0_col105[23]),
        .s(fa_s0_c105_n779_s),
        .c_out(fa_s0_c105_n779_c)
    );

    fa fa_s0_c105_n780 (
        .a(stage0_col105[24]),
        .b(stage0_col105[25]),
        .c_in(stage0_col105[26]),
        .s(fa_s0_c105_n780_s),
        .c_out(fa_s0_c105_n780_c)
    );

    fa fa_s0_c105_n781 (
        .a(stage0_col105[27]),
        .b(stage0_col105[28]),
        .c_in(stage0_col105[29]),
        .s(fa_s0_c105_n781_s),
        .c_out(fa_s0_c105_n781_c)
    );

    fa fa_s0_c106_n782 (
        .a(stage0_col106[0]),
        .b(stage0_col106[1]),
        .c_in(stage0_col106[2]),
        .s(fa_s0_c106_n782_s),
        .c_out(fa_s0_c106_n782_c)
    );

    fa fa_s0_c106_n783 (
        .a(stage0_col106[3]),
        .b(stage0_col106[4]),
        .c_in(stage0_col106[5]),
        .s(fa_s0_c106_n783_s),
        .c_out(fa_s0_c106_n783_c)
    );

    fa fa_s0_c106_n784 (
        .a(stage0_col106[6]),
        .b(stage0_col106[7]),
        .c_in(stage0_col106[8]),
        .s(fa_s0_c106_n784_s),
        .c_out(fa_s0_c106_n784_c)
    );

    fa fa_s0_c106_n785 (
        .a(stage0_col106[9]),
        .b(stage0_col106[10]),
        .c_in(stage0_col106[11]),
        .s(fa_s0_c106_n785_s),
        .c_out(fa_s0_c106_n785_c)
    );

    fa fa_s0_c106_n786 (
        .a(stage0_col106[12]),
        .b(stage0_col106[13]),
        .c_in(stage0_col106[14]),
        .s(fa_s0_c106_n786_s),
        .c_out(fa_s0_c106_n786_c)
    );

    fa fa_s0_c106_n787 (
        .a(stage0_col106[15]),
        .b(stage0_col106[16]),
        .c_in(stage0_col106[17]),
        .s(fa_s0_c106_n787_s),
        .c_out(fa_s0_c106_n787_c)
    );

    fa fa_s0_c106_n788 (
        .a(stage0_col106[18]),
        .b(stage0_col106[19]),
        .c_in(stage0_col106[20]),
        .s(fa_s0_c106_n788_s),
        .c_out(fa_s0_c106_n788_c)
    );

    fa fa_s0_c106_n789 (
        .a(stage0_col106[21]),
        .b(stage0_col106[22]),
        .c_in(stage0_col106[23]),
        .s(fa_s0_c106_n789_s),
        .c_out(fa_s0_c106_n789_c)
    );

    fa fa_s0_c106_n790 (
        .a(stage0_col106[24]),
        .b(stage0_col106[25]),
        .c_in(stage0_col106[26]),
        .s(fa_s0_c106_n790_s),
        .c_out(fa_s0_c106_n790_c)
    );

    fa fa_s0_c106_n791 (
        .a(stage0_col106[27]),
        .b(stage0_col106[28]),
        .c_in(stage0_col106[29]),
        .s(fa_s0_c106_n791_s),
        .c_out(fa_s0_c106_n791_c)
    );

    fa fa_s0_c106_n792 (
        .a(stage0_col106[30]),
        .b(stage0_col106[31]),
        .c_in(stage0_col106[32]),
        .s(fa_s0_c106_n792_s),
        .c_out(fa_s0_c106_n792_c)
    );

    fa fa_s0_c107_n793 (
        .a(stage0_col107[0]),
        .b(stage0_col107[1]),
        .c_in(stage0_col107[2]),
        .s(fa_s0_c107_n793_s),
        .c_out(fa_s0_c107_n793_c)
    );

    fa fa_s0_c107_n794 (
        .a(stage0_col107[3]),
        .b(stage0_col107[4]),
        .c_in(stage0_col107[5]),
        .s(fa_s0_c107_n794_s),
        .c_out(fa_s0_c107_n794_c)
    );

    fa fa_s0_c107_n795 (
        .a(stage0_col107[6]),
        .b(stage0_col107[7]),
        .c_in(stage0_col107[8]),
        .s(fa_s0_c107_n795_s),
        .c_out(fa_s0_c107_n795_c)
    );

    fa fa_s0_c107_n796 (
        .a(stage0_col107[9]),
        .b(stage0_col107[10]),
        .c_in(stage0_col107[11]),
        .s(fa_s0_c107_n796_s),
        .c_out(fa_s0_c107_n796_c)
    );

    fa fa_s0_c107_n797 (
        .a(stage0_col107[12]),
        .b(stage0_col107[13]),
        .c_in(stage0_col107[14]),
        .s(fa_s0_c107_n797_s),
        .c_out(fa_s0_c107_n797_c)
    );

    fa fa_s0_c107_n798 (
        .a(stage0_col107[15]),
        .b(stage0_col107[16]),
        .c_in(stage0_col107[17]),
        .s(fa_s0_c107_n798_s),
        .c_out(fa_s0_c107_n798_c)
    );

    fa fa_s0_c107_n799 (
        .a(stage0_col107[18]),
        .b(stage0_col107[19]),
        .c_in(stage0_col107[20]),
        .s(fa_s0_c107_n799_s),
        .c_out(fa_s0_c107_n799_c)
    );

    fa fa_s0_c107_n800 (
        .a(stage0_col107[21]),
        .b(stage0_col107[22]),
        .c_in(stage0_col107[23]),
        .s(fa_s0_c107_n800_s),
        .c_out(fa_s0_c107_n800_c)
    );

    fa fa_s0_c107_n801 (
        .a(stage0_col107[24]),
        .b(stage0_col107[25]),
        .c_in(stage0_col107[26]),
        .s(fa_s0_c107_n801_s),
        .c_out(fa_s0_c107_n801_c)
    );

    fa fa_s0_c107_n802 (
        .a(stage0_col107[27]),
        .b(stage0_col107[28]),
        .c_in(stage0_col107[29]),
        .s(fa_s0_c107_n802_s),
        .c_out(fa_s0_c107_n802_c)
    );

    fa fa_s0_c108_n803 (
        .a(stage0_col108[0]),
        .b(stage0_col108[1]),
        .c_in(stage0_col108[2]),
        .s(fa_s0_c108_n803_s),
        .c_out(fa_s0_c108_n803_c)
    );

    fa fa_s0_c108_n804 (
        .a(stage0_col108[3]),
        .b(stage0_col108[4]),
        .c_in(stage0_col108[5]),
        .s(fa_s0_c108_n804_s),
        .c_out(fa_s0_c108_n804_c)
    );

    fa fa_s0_c108_n805 (
        .a(stage0_col108[6]),
        .b(stage0_col108[7]),
        .c_in(stage0_col108[8]),
        .s(fa_s0_c108_n805_s),
        .c_out(fa_s0_c108_n805_c)
    );

    fa fa_s0_c108_n806 (
        .a(stage0_col108[9]),
        .b(stage0_col108[10]),
        .c_in(stage0_col108[11]),
        .s(fa_s0_c108_n806_s),
        .c_out(fa_s0_c108_n806_c)
    );

    fa fa_s0_c108_n807 (
        .a(stage0_col108[12]),
        .b(stage0_col108[13]),
        .c_in(stage0_col108[14]),
        .s(fa_s0_c108_n807_s),
        .c_out(fa_s0_c108_n807_c)
    );

    fa fa_s0_c108_n808 (
        .a(stage0_col108[15]),
        .b(stage0_col108[16]),
        .c_in(stage0_col108[17]),
        .s(fa_s0_c108_n808_s),
        .c_out(fa_s0_c108_n808_c)
    );

    fa fa_s0_c108_n809 (
        .a(stage0_col108[18]),
        .b(stage0_col108[19]),
        .c_in(stage0_col108[20]),
        .s(fa_s0_c108_n809_s),
        .c_out(fa_s0_c108_n809_c)
    );

    fa fa_s0_c108_n810 (
        .a(stage0_col108[21]),
        .b(stage0_col108[22]),
        .c_in(stage0_col108[23]),
        .s(fa_s0_c108_n810_s),
        .c_out(fa_s0_c108_n810_c)
    );

    fa fa_s0_c108_n811 (
        .a(stage0_col108[24]),
        .b(stage0_col108[25]),
        .c_in(stage0_col108[26]),
        .s(fa_s0_c108_n811_s),
        .c_out(fa_s0_c108_n811_c)
    );

    fa fa_s0_c108_n812 (
        .a(stage0_col108[27]),
        .b(stage0_col108[28]),
        .c_in(stage0_col108[29]),
        .s(fa_s0_c108_n812_s),
        .c_out(fa_s0_c108_n812_c)
    );

    fa fa_s0_c108_n813 (
        .a(stage0_col108[30]),
        .b(stage0_col108[31]),
        .c_in(stage0_col108[32]),
        .s(fa_s0_c108_n813_s),
        .c_out(fa_s0_c108_n813_c)
    );

    fa fa_s0_c109_n814 (
        .a(stage0_col109[0]),
        .b(stage0_col109[1]),
        .c_in(stage0_col109[2]),
        .s(fa_s0_c109_n814_s),
        .c_out(fa_s0_c109_n814_c)
    );

    fa fa_s0_c109_n815 (
        .a(stage0_col109[3]),
        .b(stage0_col109[4]),
        .c_in(stage0_col109[5]),
        .s(fa_s0_c109_n815_s),
        .c_out(fa_s0_c109_n815_c)
    );

    fa fa_s0_c109_n816 (
        .a(stage0_col109[6]),
        .b(stage0_col109[7]),
        .c_in(stage0_col109[8]),
        .s(fa_s0_c109_n816_s),
        .c_out(fa_s0_c109_n816_c)
    );

    fa fa_s0_c109_n817 (
        .a(stage0_col109[9]),
        .b(stage0_col109[10]),
        .c_in(stage0_col109[11]),
        .s(fa_s0_c109_n817_s),
        .c_out(fa_s0_c109_n817_c)
    );

    fa fa_s0_c109_n818 (
        .a(stage0_col109[12]),
        .b(stage0_col109[13]),
        .c_in(stage0_col109[14]),
        .s(fa_s0_c109_n818_s),
        .c_out(fa_s0_c109_n818_c)
    );

    fa fa_s0_c109_n819 (
        .a(stage0_col109[15]),
        .b(stage0_col109[16]),
        .c_in(stage0_col109[17]),
        .s(fa_s0_c109_n819_s),
        .c_out(fa_s0_c109_n819_c)
    );

    fa fa_s0_c109_n820 (
        .a(stage0_col109[18]),
        .b(stage0_col109[19]),
        .c_in(stage0_col109[20]),
        .s(fa_s0_c109_n820_s),
        .c_out(fa_s0_c109_n820_c)
    );

    fa fa_s0_c109_n821 (
        .a(stage0_col109[21]),
        .b(stage0_col109[22]),
        .c_in(stage0_col109[23]),
        .s(fa_s0_c109_n821_s),
        .c_out(fa_s0_c109_n821_c)
    );

    fa fa_s0_c109_n822 (
        .a(stage0_col109[24]),
        .b(stage0_col109[25]),
        .c_in(stage0_col109[26]),
        .s(fa_s0_c109_n822_s),
        .c_out(fa_s0_c109_n822_c)
    );

    fa fa_s0_c109_n823 (
        .a(stage0_col109[27]),
        .b(stage0_col109[28]),
        .c_in(stage0_col109[29]),
        .s(fa_s0_c109_n823_s),
        .c_out(fa_s0_c109_n823_c)
    );

    fa fa_s0_c110_n824 (
        .a(stage0_col110[0]),
        .b(stage0_col110[1]),
        .c_in(stage0_col110[2]),
        .s(fa_s0_c110_n824_s),
        .c_out(fa_s0_c110_n824_c)
    );

    fa fa_s0_c110_n825 (
        .a(stage0_col110[3]),
        .b(stage0_col110[4]),
        .c_in(stage0_col110[5]),
        .s(fa_s0_c110_n825_s),
        .c_out(fa_s0_c110_n825_c)
    );

    fa fa_s0_c110_n826 (
        .a(stage0_col110[6]),
        .b(stage0_col110[7]),
        .c_in(stage0_col110[8]),
        .s(fa_s0_c110_n826_s),
        .c_out(fa_s0_c110_n826_c)
    );

    fa fa_s0_c110_n827 (
        .a(stage0_col110[9]),
        .b(stage0_col110[10]),
        .c_in(stage0_col110[11]),
        .s(fa_s0_c110_n827_s),
        .c_out(fa_s0_c110_n827_c)
    );

    fa fa_s0_c110_n828 (
        .a(stage0_col110[12]),
        .b(stage0_col110[13]),
        .c_in(stage0_col110[14]),
        .s(fa_s0_c110_n828_s),
        .c_out(fa_s0_c110_n828_c)
    );

    fa fa_s0_c110_n829 (
        .a(stage0_col110[15]),
        .b(stage0_col110[16]),
        .c_in(stage0_col110[17]),
        .s(fa_s0_c110_n829_s),
        .c_out(fa_s0_c110_n829_c)
    );

    fa fa_s0_c110_n830 (
        .a(stage0_col110[18]),
        .b(stage0_col110[19]),
        .c_in(stage0_col110[20]),
        .s(fa_s0_c110_n830_s),
        .c_out(fa_s0_c110_n830_c)
    );

    fa fa_s0_c110_n831 (
        .a(stage0_col110[21]),
        .b(stage0_col110[22]),
        .c_in(stage0_col110[23]),
        .s(fa_s0_c110_n831_s),
        .c_out(fa_s0_c110_n831_c)
    );

    fa fa_s0_c110_n832 (
        .a(stage0_col110[24]),
        .b(stage0_col110[25]),
        .c_in(stage0_col110[26]),
        .s(fa_s0_c110_n832_s),
        .c_out(fa_s0_c110_n832_c)
    );

    fa fa_s0_c110_n833 (
        .a(stage0_col110[27]),
        .b(stage0_col110[28]),
        .c_in(stage0_col110[29]),
        .s(fa_s0_c110_n833_s),
        .c_out(fa_s0_c110_n833_c)
    );

    fa fa_s0_c110_n834 (
        .a(stage0_col110[30]),
        .b(stage0_col110[31]),
        .c_in(stage0_col110[32]),
        .s(fa_s0_c110_n834_s),
        .c_out(fa_s0_c110_n834_c)
    );

    fa fa_s0_c111_n835 (
        .a(stage0_col111[0]),
        .b(stage0_col111[1]),
        .c_in(stage0_col111[2]),
        .s(fa_s0_c111_n835_s),
        .c_out(fa_s0_c111_n835_c)
    );

    fa fa_s0_c111_n836 (
        .a(stage0_col111[3]),
        .b(stage0_col111[4]),
        .c_in(stage0_col111[5]),
        .s(fa_s0_c111_n836_s),
        .c_out(fa_s0_c111_n836_c)
    );

    fa fa_s0_c111_n837 (
        .a(stage0_col111[6]),
        .b(stage0_col111[7]),
        .c_in(stage0_col111[8]),
        .s(fa_s0_c111_n837_s),
        .c_out(fa_s0_c111_n837_c)
    );

    fa fa_s0_c111_n838 (
        .a(stage0_col111[9]),
        .b(stage0_col111[10]),
        .c_in(stage0_col111[11]),
        .s(fa_s0_c111_n838_s),
        .c_out(fa_s0_c111_n838_c)
    );

    fa fa_s0_c111_n839 (
        .a(stage0_col111[12]),
        .b(stage0_col111[13]),
        .c_in(stage0_col111[14]),
        .s(fa_s0_c111_n839_s),
        .c_out(fa_s0_c111_n839_c)
    );

    fa fa_s0_c111_n840 (
        .a(stage0_col111[15]),
        .b(stage0_col111[16]),
        .c_in(stage0_col111[17]),
        .s(fa_s0_c111_n840_s),
        .c_out(fa_s0_c111_n840_c)
    );

    fa fa_s0_c111_n841 (
        .a(stage0_col111[18]),
        .b(stage0_col111[19]),
        .c_in(stage0_col111[20]),
        .s(fa_s0_c111_n841_s),
        .c_out(fa_s0_c111_n841_c)
    );

    fa fa_s0_c111_n842 (
        .a(stage0_col111[21]),
        .b(stage0_col111[22]),
        .c_in(stage0_col111[23]),
        .s(fa_s0_c111_n842_s),
        .c_out(fa_s0_c111_n842_c)
    );

    fa fa_s0_c111_n843 (
        .a(stage0_col111[24]),
        .b(stage0_col111[25]),
        .c_in(stage0_col111[26]),
        .s(fa_s0_c111_n843_s),
        .c_out(fa_s0_c111_n843_c)
    );

    fa fa_s0_c111_n844 (
        .a(stage0_col111[27]),
        .b(stage0_col111[28]),
        .c_in(stage0_col111[29]),
        .s(fa_s0_c111_n844_s),
        .c_out(fa_s0_c111_n844_c)
    );

    fa fa_s0_c112_n845 (
        .a(stage0_col112[0]),
        .b(stage0_col112[1]),
        .c_in(stage0_col112[2]),
        .s(fa_s0_c112_n845_s),
        .c_out(fa_s0_c112_n845_c)
    );

    fa fa_s0_c112_n846 (
        .a(stage0_col112[3]),
        .b(stage0_col112[4]),
        .c_in(stage0_col112[5]),
        .s(fa_s0_c112_n846_s),
        .c_out(fa_s0_c112_n846_c)
    );

    fa fa_s0_c112_n847 (
        .a(stage0_col112[6]),
        .b(stage0_col112[7]),
        .c_in(stage0_col112[8]),
        .s(fa_s0_c112_n847_s),
        .c_out(fa_s0_c112_n847_c)
    );

    fa fa_s0_c112_n848 (
        .a(stage0_col112[9]),
        .b(stage0_col112[10]),
        .c_in(stage0_col112[11]),
        .s(fa_s0_c112_n848_s),
        .c_out(fa_s0_c112_n848_c)
    );

    fa fa_s0_c112_n849 (
        .a(stage0_col112[12]),
        .b(stage0_col112[13]),
        .c_in(stage0_col112[14]),
        .s(fa_s0_c112_n849_s),
        .c_out(fa_s0_c112_n849_c)
    );

    fa fa_s0_c112_n850 (
        .a(stage0_col112[15]),
        .b(stage0_col112[16]),
        .c_in(stage0_col112[17]),
        .s(fa_s0_c112_n850_s),
        .c_out(fa_s0_c112_n850_c)
    );

    fa fa_s0_c112_n851 (
        .a(stage0_col112[18]),
        .b(stage0_col112[19]),
        .c_in(stage0_col112[20]),
        .s(fa_s0_c112_n851_s),
        .c_out(fa_s0_c112_n851_c)
    );

    fa fa_s0_c112_n852 (
        .a(stage0_col112[21]),
        .b(stage0_col112[22]),
        .c_in(stage0_col112[23]),
        .s(fa_s0_c112_n852_s),
        .c_out(fa_s0_c112_n852_c)
    );

    fa fa_s0_c112_n853 (
        .a(stage0_col112[24]),
        .b(stage0_col112[25]),
        .c_in(stage0_col112[26]),
        .s(fa_s0_c112_n853_s),
        .c_out(fa_s0_c112_n853_c)
    );

    fa fa_s0_c112_n854 (
        .a(stage0_col112[27]),
        .b(stage0_col112[28]),
        .c_in(stage0_col112[29]),
        .s(fa_s0_c112_n854_s),
        .c_out(fa_s0_c112_n854_c)
    );

    fa fa_s0_c112_n855 (
        .a(stage0_col112[30]),
        .b(stage0_col112[31]),
        .c_in(stage0_col112[32]),
        .s(fa_s0_c112_n855_s),
        .c_out(fa_s0_c112_n855_c)
    );

    fa fa_s0_c113_n856 (
        .a(stage0_col113[0]),
        .b(stage0_col113[1]),
        .c_in(stage0_col113[2]),
        .s(fa_s0_c113_n856_s),
        .c_out(fa_s0_c113_n856_c)
    );

    fa fa_s0_c113_n857 (
        .a(stage0_col113[3]),
        .b(stage0_col113[4]),
        .c_in(stage0_col113[5]),
        .s(fa_s0_c113_n857_s),
        .c_out(fa_s0_c113_n857_c)
    );

    fa fa_s0_c113_n858 (
        .a(stage0_col113[6]),
        .b(stage0_col113[7]),
        .c_in(stage0_col113[8]),
        .s(fa_s0_c113_n858_s),
        .c_out(fa_s0_c113_n858_c)
    );

    fa fa_s0_c113_n859 (
        .a(stage0_col113[9]),
        .b(stage0_col113[10]),
        .c_in(stage0_col113[11]),
        .s(fa_s0_c113_n859_s),
        .c_out(fa_s0_c113_n859_c)
    );

    fa fa_s0_c113_n860 (
        .a(stage0_col113[12]),
        .b(stage0_col113[13]),
        .c_in(stage0_col113[14]),
        .s(fa_s0_c113_n860_s),
        .c_out(fa_s0_c113_n860_c)
    );

    fa fa_s0_c113_n861 (
        .a(stage0_col113[15]),
        .b(stage0_col113[16]),
        .c_in(stage0_col113[17]),
        .s(fa_s0_c113_n861_s),
        .c_out(fa_s0_c113_n861_c)
    );

    fa fa_s0_c113_n862 (
        .a(stage0_col113[18]),
        .b(stage0_col113[19]),
        .c_in(stage0_col113[20]),
        .s(fa_s0_c113_n862_s),
        .c_out(fa_s0_c113_n862_c)
    );

    fa fa_s0_c113_n863 (
        .a(stage0_col113[21]),
        .b(stage0_col113[22]),
        .c_in(stage0_col113[23]),
        .s(fa_s0_c113_n863_s),
        .c_out(fa_s0_c113_n863_c)
    );

    fa fa_s0_c113_n864 (
        .a(stage0_col113[24]),
        .b(stage0_col113[25]),
        .c_in(stage0_col113[26]),
        .s(fa_s0_c113_n864_s),
        .c_out(fa_s0_c113_n864_c)
    );

    fa fa_s0_c113_n865 (
        .a(stage0_col113[27]),
        .b(stage0_col113[28]),
        .c_in(stage0_col113[29]),
        .s(fa_s0_c113_n865_s),
        .c_out(fa_s0_c113_n865_c)
    );

    fa fa_s0_c114_n866 (
        .a(stage0_col114[0]),
        .b(stage0_col114[1]),
        .c_in(stage0_col114[2]),
        .s(fa_s0_c114_n866_s),
        .c_out(fa_s0_c114_n866_c)
    );

    fa fa_s0_c114_n867 (
        .a(stage0_col114[3]),
        .b(stage0_col114[4]),
        .c_in(stage0_col114[5]),
        .s(fa_s0_c114_n867_s),
        .c_out(fa_s0_c114_n867_c)
    );

    fa fa_s0_c114_n868 (
        .a(stage0_col114[6]),
        .b(stage0_col114[7]),
        .c_in(stage0_col114[8]),
        .s(fa_s0_c114_n868_s),
        .c_out(fa_s0_c114_n868_c)
    );

    fa fa_s0_c114_n869 (
        .a(stage0_col114[9]),
        .b(stage0_col114[10]),
        .c_in(stage0_col114[11]),
        .s(fa_s0_c114_n869_s),
        .c_out(fa_s0_c114_n869_c)
    );

    fa fa_s0_c114_n870 (
        .a(stage0_col114[12]),
        .b(stage0_col114[13]),
        .c_in(stage0_col114[14]),
        .s(fa_s0_c114_n870_s),
        .c_out(fa_s0_c114_n870_c)
    );

    fa fa_s0_c114_n871 (
        .a(stage0_col114[15]),
        .b(stage0_col114[16]),
        .c_in(stage0_col114[17]),
        .s(fa_s0_c114_n871_s),
        .c_out(fa_s0_c114_n871_c)
    );

    fa fa_s0_c114_n872 (
        .a(stage0_col114[18]),
        .b(stage0_col114[19]),
        .c_in(stage0_col114[20]),
        .s(fa_s0_c114_n872_s),
        .c_out(fa_s0_c114_n872_c)
    );

    fa fa_s0_c114_n873 (
        .a(stage0_col114[21]),
        .b(stage0_col114[22]),
        .c_in(stage0_col114[23]),
        .s(fa_s0_c114_n873_s),
        .c_out(fa_s0_c114_n873_c)
    );

    fa fa_s0_c114_n874 (
        .a(stage0_col114[24]),
        .b(stage0_col114[25]),
        .c_in(stage0_col114[26]),
        .s(fa_s0_c114_n874_s),
        .c_out(fa_s0_c114_n874_c)
    );

    fa fa_s0_c114_n875 (
        .a(stage0_col114[27]),
        .b(stage0_col114[28]),
        .c_in(stage0_col114[29]),
        .s(fa_s0_c114_n875_s),
        .c_out(fa_s0_c114_n875_c)
    );

    fa fa_s0_c114_n876 (
        .a(stage0_col114[30]),
        .b(stage0_col114[31]),
        .c_in(stage0_col114[32]),
        .s(fa_s0_c114_n876_s),
        .c_out(fa_s0_c114_n876_c)
    );

    fa fa_s0_c115_n877 (
        .a(stage0_col115[0]),
        .b(stage0_col115[1]),
        .c_in(stage0_col115[2]),
        .s(fa_s0_c115_n877_s),
        .c_out(fa_s0_c115_n877_c)
    );

    fa fa_s0_c115_n878 (
        .a(stage0_col115[3]),
        .b(stage0_col115[4]),
        .c_in(stage0_col115[5]),
        .s(fa_s0_c115_n878_s),
        .c_out(fa_s0_c115_n878_c)
    );

    fa fa_s0_c115_n879 (
        .a(stage0_col115[6]),
        .b(stage0_col115[7]),
        .c_in(stage0_col115[8]),
        .s(fa_s0_c115_n879_s),
        .c_out(fa_s0_c115_n879_c)
    );

    fa fa_s0_c115_n880 (
        .a(stage0_col115[9]),
        .b(stage0_col115[10]),
        .c_in(stage0_col115[11]),
        .s(fa_s0_c115_n880_s),
        .c_out(fa_s0_c115_n880_c)
    );

    fa fa_s0_c115_n881 (
        .a(stage0_col115[12]),
        .b(stage0_col115[13]),
        .c_in(stage0_col115[14]),
        .s(fa_s0_c115_n881_s),
        .c_out(fa_s0_c115_n881_c)
    );

    fa fa_s0_c115_n882 (
        .a(stage0_col115[15]),
        .b(stage0_col115[16]),
        .c_in(stage0_col115[17]),
        .s(fa_s0_c115_n882_s),
        .c_out(fa_s0_c115_n882_c)
    );

    fa fa_s0_c115_n883 (
        .a(stage0_col115[18]),
        .b(stage0_col115[19]),
        .c_in(stage0_col115[20]),
        .s(fa_s0_c115_n883_s),
        .c_out(fa_s0_c115_n883_c)
    );

    fa fa_s0_c115_n884 (
        .a(stage0_col115[21]),
        .b(stage0_col115[22]),
        .c_in(stage0_col115[23]),
        .s(fa_s0_c115_n884_s),
        .c_out(fa_s0_c115_n884_c)
    );

    fa fa_s0_c115_n885 (
        .a(stage0_col115[24]),
        .b(stage0_col115[25]),
        .c_in(stage0_col115[26]),
        .s(fa_s0_c115_n885_s),
        .c_out(fa_s0_c115_n885_c)
    );

    fa fa_s0_c115_n886 (
        .a(stage0_col115[27]),
        .b(stage0_col115[28]),
        .c_in(stage0_col115[29]),
        .s(fa_s0_c115_n886_s),
        .c_out(fa_s0_c115_n886_c)
    );

    fa fa_s0_c116_n887 (
        .a(stage0_col116[0]),
        .b(stage0_col116[1]),
        .c_in(stage0_col116[2]),
        .s(fa_s0_c116_n887_s),
        .c_out(fa_s0_c116_n887_c)
    );

    fa fa_s0_c116_n888 (
        .a(stage0_col116[3]),
        .b(stage0_col116[4]),
        .c_in(stage0_col116[5]),
        .s(fa_s0_c116_n888_s),
        .c_out(fa_s0_c116_n888_c)
    );

    fa fa_s0_c116_n889 (
        .a(stage0_col116[6]),
        .b(stage0_col116[7]),
        .c_in(stage0_col116[8]),
        .s(fa_s0_c116_n889_s),
        .c_out(fa_s0_c116_n889_c)
    );

    fa fa_s0_c116_n890 (
        .a(stage0_col116[9]),
        .b(stage0_col116[10]),
        .c_in(stage0_col116[11]),
        .s(fa_s0_c116_n890_s),
        .c_out(fa_s0_c116_n890_c)
    );

    fa fa_s0_c116_n891 (
        .a(stage0_col116[12]),
        .b(stage0_col116[13]),
        .c_in(stage0_col116[14]),
        .s(fa_s0_c116_n891_s),
        .c_out(fa_s0_c116_n891_c)
    );

    fa fa_s0_c116_n892 (
        .a(stage0_col116[15]),
        .b(stage0_col116[16]),
        .c_in(stage0_col116[17]),
        .s(fa_s0_c116_n892_s),
        .c_out(fa_s0_c116_n892_c)
    );

    fa fa_s0_c116_n893 (
        .a(stage0_col116[18]),
        .b(stage0_col116[19]),
        .c_in(stage0_col116[20]),
        .s(fa_s0_c116_n893_s),
        .c_out(fa_s0_c116_n893_c)
    );

    fa fa_s0_c116_n894 (
        .a(stage0_col116[21]),
        .b(stage0_col116[22]),
        .c_in(stage0_col116[23]),
        .s(fa_s0_c116_n894_s),
        .c_out(fa_s0_c116_n894_c)
    );

    fa fa_s0_c116_n895 (
        .a(stage0_col116[24]),
        .b(stage0_col116[25]),
        .c_in(stage0_col116[26]),
        .s(fa_s0_c116_n895_s),
        .c_out(fa_s0_c116_n895_c)
    );

    fa fa_s0_c116_n896 (
        .a(stage0_col116[27]),
        .b(stage0_col116[28]),
        .c_in(stage0_col116[29]),
        .s(fa_s0_c116_n896_s),
        .c_out(fa_s0_c116_n896_c)
    );

    fa fa_s0_c116_n897 (
        .a(stage0_col116[30]),
        .b(stage0_col116[31]),
        .c_in(stage0_col116[32]),
        .s(fa_s0_c116_n897_s),
        .c_out(fa_s0_c116_n897_c)
    );

    fa fa_s0_c117_n898 (
        .a(stage0_col117[0]),
        .b(stage0_col117[1]),
        .c_in(stage0_col117[2]),
        .s(fa_s0_c117_n898_s),
        .c_out(fa_s0_c117_n898_c)
    );

    fa fa_s0_c117_n899 (
        .a(stage0_col117[3]),
        .b(stage0_col117[4]),
        .c_in(stage0_col117[5]),
        .s(fa_s0_c117_n899_s),
        .c_out(fa_s0_c117_n899_c)
    );

    fa fa_s0_c117_n900 (
        .a(stage0_col117[6]),
        .b(stage0_col117[7]),
        .c_in(stage0_col117[8]),
        .s(fa_s0_c117_n900_s),
        .c_out(fa_s0_c117_n900_c)
    );

    fa fa_s0_c117_n901 (
        .a(stage0_col117[9]),
        .b(stage0_col117[10]),
        .c_in(stage0_col117[11]),
        .s(fa_s0_c117_n901_s),
        .c_out(fa_s0_c117_n901_c)
    );

    fa fa_s0_c117_n902 (
        .a(stage0_col117[12]),
        .b(stage0_col117[13]),
        .c_in(stage0_col117[14]),
        .s(fa_s0_c117_n902_s),
        .c_out(fa_s0_c117_n902_c)
    );

    fa fa_s0_c117_n903 (
        .a(stage0_col117[15]),
        .b(stage0_col117[16]),
        .c_in(stage0_col117[17]),
        .s(fa_s0_c117_n903_s),
        .c_out(fa_s0_c117_n903_c)
    );

    fa fa_s0_c117_n904 (
        .a(stage0_col117[18]),
        .b(stage0_col117[19]),
        .c_in(stage0_col117[20]),
        .s(fa_s0_c117_n904_s),
        .c_out(fa_s0_c117_n904_c)
    );

    fa fa_s0_c117_n905 (
        .a(stage0_col117[21]),
        .b(stage0_col117[22]),
        .c_in(stage0_col117[23]),
        .s(fa_s0_c117_n905_s),
        .c_out(fa_s0_c117_n905_c)
    );

    fa fa_s0_c117_n906 (
        .a(stage0_col117[24]),
        .b(stage0_col117[25]),
        .c_in(stage0_col117[26]),
        .s(fa_s0_c117_n906_s),
        .c_out(fa_s0_c117_n906_c)
    );

    fa fa_s0_c117_n907 (
        .a(stage0_col117[27]),
        .b(stage0_col117[28]),
        .c_in(stage0_col117[29]),
        .s(fa_s0_c117_n907_s),
        .c_out(fa_s0_c117_n907_c)
    );

    fa fa_s0_c118_n908 (
        .a(stage0_col118[0]),
        .b(stage0_col118[1]),
        .c_in(stage0_col118[2]),
        .s(fa_s0_c118_n908_s),
        .c_out(fa_s0_c118_n908_c)
    );

    fa fa_s0_c118_n909 (
        .a(stage0_col118[3]),
        .b(stage0_col118[4]),
        .c_in(stage0_col118[5]),
        .s(fa_s0_c118_n909_s),
        .c_out(fa_s0_c118_n909_c)
    );

    fa fa_s0_c118_n910 (
        .a(stage0_col118[6]),
        .b(stage0_col118[7]),
        .c_in(stage0_col118[8]),
        .s(fa_s0_c118_n910_s),
        .c_out(fa_s0_c118_n910_c)
    );

    fa fa_s0_c118_n911 (
        .a(stage0_col118[9]),
        .b(stage0_col118[10]),
        .c_in(stage0_col118[11]),
        .s(fa_s0_c118_n911_s),
        .c_out(fa_s0_c118_n911_c)
    );

    fa fa_s0_c118_n912 (
        .a(stage0_col118[12]),
        .b(stage0_col118[13]),
        .c_in(stage0_col118[14]),
        .s(fa_s0_c118_n912_s),
        .c_out(fa_s0_c118_n912_c)
    );

    fa fa_s0_c118_n913 (
        .a(stage0_col118[15]),
        .b(stage0_col118[16]),
        .c_in(stage0_col118[17]),
        .s(fa_s0_c118_n913_s),
        .c_out(fa_s0_c118_n913_c)
    );

    fa fa_s0_c118_n914 (
        .a(stage0_col118[18]),
        .b(stage0_col118[19]),
        .c_in(stage0_col118[20]),
        .s(fa_s0_c118_n914_s),
        .c_out(fa_s0_c118_n914_c)
    );

    fa fa_s0_c118_n915 (
        .a(stage0_col118[21]),
        .b(stage0_col118[22]),
        .c_in(stage0_col118[23]),
        .s(fa_s0_c118_n915_s),
        .c_out(fa_s0_c118_n915_c)
    );

    fa fa_s0_c118_n916 (
        .a(stage0_col118[24]),
        .b(stage0_col118[25]),
        .c_in(stage0_col118[26]),
        .s(fa_s0_c118_n916_s),
        .c_out(fa_s0_c118_n916_c)
    );

    fa fa_s0_c118_n917 (
        .a(stage0_col118[27]),
        .b(stage0_col118[28]),
        .c_in(stage0_col118[29]),
        .s(fa_s0_c118_n917_s),
        .c_out(fa_s0_c118_n917_c)
    );

    fa fa_s0_c118_n918 (
        .a(stage0_col118[30]),
        .b(stage0_col118[31]),
        .c_in(stage0_col118[32]),
        .s(fa_s0_c118_n918_s),
        .c_out(fa_s0_c118_n918_c)
    );

    fa fa_s0_c119_n919 (
        .a(stage0_col119[0]),
        .b(stage0_col119[1]),
        .c_in(stage0_col119[2]),
        .s(fa_s0_c119_n919_s),
        .c_out(fa_s0_c119_n919_c)
    );

    fa fa_s0_c119_n920 (
        .a(stage0_col119[3]),
        .b(stage0_col119[4]),
        .c_in(stage0_col119[5]),
        .s(fa_s0_c119_n920_s),
        .c_out(fa_s0_c119_n920_c)
    );

    fa fa_s0_c119_n921 (
        .a(stage0_col119[6]),
        .b(stage0_col119[7]),
        .c_in(stage0_col119[8]),
        .s(fa_s0_c119_n921_s),
        .c_out(fa_s0_c119_n921_c)
    );

    fa fa_s0_c119_n922 (
        .a(stage0_col119[9]),
        .b(stage0_col119[10]),
        .c_in(stage0_col119[11]),
        .s(fa_s0_c119_n922_s),
        .c_out(fa_s0_c119_n922_c)
    );

    fa fa_s0_c119_n923 (
        .a(stage0_col119[12]),
        .b(stage0_col119[13]),
        .c_in(stage0_col119[14]),
        .s(fa_s0_c119_n923_s),
        .c_out(fa_s0_c119_n923_c)
    );

    fa fa_s0_c119_n924 (
        .a(stage0_col119[15]),
        .b(stage0_col119[16]),
        .c_in(stage0_col119[17]),
        .s(fa_s0_c119_n924_s),
        .c_out(fa_s0_c119_n924_c)
    );

    fa fa_s0_c119_n925 (
        .a(stage0_col119[18]),
        .b(stage0_col119[19]),
        .c_in(stage0_col119[20]),
        .s(fa_s0_c119_n925_s),
        .c_out(fa_s0_c119_n925_c)
    );

    fa fa_s0_c119_n926 (
        .a(stage0_col119[21]),
        .b(stage0_col119[22]),
        .c_in(stage0_col119[23]),
        .s(fa_s0_c119_n926_s),
        .c_out(fa_s0_c119_n926_c)
    );

    fa fa_s0_c119_n927 (
        .a(stage0_col119[24]),
        .b(stage0_col119[25]),
        .c_in(stage0_col119[26]),
        .s(fa_s0_c119_n927_s),
        .c_out(fa_s0_c119_n927_c)
    );

    fa fa_s0_c119_n928 (
        .a(stage0_col119[27]),
        .b(stage0_col119[28]),
        .c_in(stage0_col119[29]),
        .s(fa_s0_c119_n928_s),
        .c_out(fa_s0_c119_n928_c)
    );

    fa fa_s0_c120_n929 (
        .a(stage0_col120[0]),
        .b(stage0_col120[1]),
        .c_in(stage0_col120[2]),
        .s(fa_s0_c120_n929_s),
        .c_out(fa_s0_c120_n929_c)
    );

    fa fa_s0_c120_n930 (
        .a(stage0_col120[3]),
        .b(stage0_col120[4]),
        .c_in(stage0_col120[5]),
        .s(fa_s0_c120_n930_s),
        .c_out(fa_s0_c120_n930_c)
    );

    fa fa_s0_c120_n931 (
        .a(stage0_col120[6]),
        .b(stage0_col120[7]),
        .c_in(stage0_col120[8]),
        .s(fa_s0_c120_n931_s),
        .c_out(fa_s0_c120_n931_c)
    );

    fa fa_s0_c120_n932 (
        .a(stage0_col120[9]),
        .b(stage0_col120[10]),
        .c_in(stage0_col120[11]),
        .s(fa_s0_c120_n932_s),
        .c_out(fa_s0_c120_n932_c)
    );

    fa fa_s0_c120_n933 (
        .a(stage0_col120[12]),
        .b(stage0_col120[13]),
        .c_in(stage0_col120[14]),
        .s(fa_s0_c120_n933_s),
        .c_out(fa_s0_c120_n933_c)
    );

    fa fa_s0_c120_n934 (
        .a(stage0_col120[15]),
        .b(stage0_col120[16]),
        .c_in(stage0_col120[17]),
        .s(fa_s0_c120_n934_s),
        .c_out(fa_s0_c120_n934_c)
    );

    fa fa_s0_c120_n935 (
        .a(stage0_col120[18]),
        .b(stage0_col120[19]),
        .c_in(stage0_col120[20]),
        .s(fa_s0_c120_n935_s),
        .c_out(fa_s0_c120_n935_c)
    );

    fa fa_s0_c120_n936 (
        .a(stage0_col120[21]),
        .b(stage0_col120[22]),
        .c_in(stage0_col120[23]),
        .s(fa_s0_c120_n936_s),
        .c_out(fa_s0_c120_n936_c)
    );

    fa fa_s0_c120_n937 (
        .a(stage0_col120[24]),
        .b(stage0_col120[25]),
        .c_in(stage0_col120[26]),
        .s(fa_s0_c120_n937_s),
        .c_out(fa_s0_c120_n937_c)
    );

    fa fa_s0_c120_n938 (
        .a(stage0_col120[27]),
        .b(stage0_col120[28]),
        .c_in(stage0_col120[29]),
        .s(fa_s0_c120_n938_s),
        .c_out(fa_s0_c120_n938_c)
    );

    fa fa_s0_c120_n939 (
        .a(stage0_col120[30]),
        .b(stage0_col120[31]),
        .c_in(stage0_col120[32]),
        .s(fa_s0_c120_n939_s),
        .c_out(fa_s0_c120_n939_c)
    );

    fa fa_s0_c121_n940 (
        .a(stage0_col121[0]),
        .b(stage0_col121[1]),
        .c_in(stage0_col121[2]),
        .s(fa_s0_c121_n940_s),
        .c_out(fa_s0_c121_n940_c)
    );

    fa fa_s0_c121_n941 (
        .a(stage0_col121[3]),
        .b(stage0_col121[4]),
        .c_in(stage0_col121[5]),
        .s(fa_s0_c121_n941_s),
        .c_out(fa_s0_c121_n941_c)
    );

    fa fa_s0_c121_n942 (
        .a(stage0_col121[6]),
        .b(stage0_col121[7]),
        .c_in(stage0_col121[8]),
        .s(fa_s0_c121_n942_s),
        .c_out(fa_s0_c121_n942_c)
    );

    fa fa_s0_c121_n943 (
        .a(stage0_col121[9]),
        .b(stage0_col121[10]),
        .c_in(stage0_col121[11]),
        .s(fa_s0_c121_n943_s),
        .c_out(fa_s0_c121_n943_c)
    );

    fa fa_s0_c121_n944 (
        .a(stage0_col121[12]),
        .b(stage0_col121[13]),
        .c_in(stage0_col121[14]),
        .s(fa_s0_c121_n944_s),
        .c_out(fa_s0_c121_n944_c)
    );

    fa fa_s0_c121_n945 (
        .a(stage0_col121[15]),
        .b(stage0_col121[16]),
        .c_in(stage0_col121[17]),
        .s(fa_s0_c121_n945_s),
        .c_out(fa_s0_c121_n945_c)
    );

    fa fa_s0_c121_n946 (
        .a(stage0_col121[18]),
        .b(stage0_col121[19]),
        .c_in(stage0_col121[20]),
        .s(fa_s0_c121_n946_s),
        .c_out(fa_s0_c121_n946_c)
    );

    fa fa_s0_c121_n947 (
        .a(stage0_col121[21]),
        .b(stage0_col121[22]),
        .c_in(stage0_col121[23]),
        .s(fa_s0_c121_n947_s),
        .c_out(fa_s0_c121_n947_c)
    );

    fa fa_s0_c121_n948 (
        .a(stage0_col121[24]),
        .b(stage0_col121[25]),
        .c_in(stage0_col121[26]),
        .s(fa_s0_c121_n948_s),
        .c_out(fa_s0_c121_n948_c)
    );

    fa fa_s0_c121_n949 (
        .a(stage0_col121[27]),
        .b(stage0_col121[28]),
        .c_in(stage0_col121[29]),
        .s(fa_s0_c121_n949_s),
        .c_out(fa_s0_c121_n949_c)
    );

    fa fa_s0_c122_n950 (
        .a(stage0_col122[0]),
        .b(stage0_col122[1]),
        .c_in(stage0_col122[2]),
        .s(fa_s0_c122_n950_s),
        .c_out(fa_s0_c122_n950_c)
    );

    fa fa_s0_c122_n951 (
        .a(stage0_col122[3]),
        .b(stage0_col122[4]),
        .c_in(stage0_col122[5]),
        .s(fa_s0_c122_n951_s),
        .c_out(fa_s0_c122_n951_c)
    );

    fa fa_s0_c122_n952 (
        .a(stage0_col122[6]),
        .b(stage0_col122[7]),
        .c_in(stage0_col122[8]),
        .s(fa_s0_c122_n952_s),
        .c_out(fa_s0_c122_n952_c)
    );

    fa fa_s0_c122_n953 (
        .a(stage0_col122[9]),
        .b(stage0_col122[10]),
        .c_in(stage0_col122[11]),
        .s(fa_s0_c122_n953_s),
        .c_out(fa_s0_c122_n953_c)
    );

    fa fa_s0_c122_n954 (
        .a(stage0_col122[12]),
        .b(stage0_col122[13]),
        .c_in(stage0_col122[14]),
        .s(fa_s0_c122_n954_s),
        .c_out(fa_s0_c122_n954_c)
    );

    fa fa_s0_c122_n955 (
        .a(stage0_col122[15]),
        .b(stage0_col122[16]),
        .c_in(stage0_col122[17]),
        .s(fa_s0_c122_n955_s),
        .c_out(fa_s0_c122_n955_c)
    );

    fa fa_s0_c122_n956 (
        .a(stage0_col122[18]),
        .b(stage0_col122[19]),
        .c_in(stage0_col122[20]),
        .s(fa_s0_c122_n956_s),
        .c_out(fa_s0_c122_n956_c)
    );

    fa fa_s0_c122_n957 (
        .a(stage0_col122[21]),
        .b(stage0_col122[22]),
        .c_in(stage0_col122[23]),
        .s(fa_s0_c122_n957_s),
        .c_out(fa_s0_c122_n957_c)
    );

    fa fa_s0_c122_n958 (
        .a(stage0_col122[24]),
        .b(stage0_col122[25]),
        .c_in(stage0_col122[26]),
        .s(fa_s0_c122_n958_s),
        .c_out(fa_s0_c122_n958_c)
    );

    fa fa_s0_c122_n959 (
        .a(stage0_col122[27]),
        .b(stage0_col122[28]),
        .c_in(stage0_col122[29]),
        .s(fa_s0_c122_n959_s),
        .c_out(fa_s0_c122_n959_c)
    );

    fa fa_s0_c122_n960 (
        .a(stage0_col122[30]),
        .b(stage0_col122[31]),
        .c_in(stage0_col122[32]),
        .s(fa_s0_c122_n960_s),
        .c_out(fa_s0_c122_n960_c)
    );

    fa fa_s0_c123_n961 (
        .a(stage0_col123[0]),
        .b(stage0_col123[1]),
        .c_in(stage0_col123[2]),
        .s(fa_s0_c123_n961_s),
        .c_out(fa_s0_c123_n961_c)
    );

    fa fa_s0_c123_n962 (
        .a(stage0_col123[3]),
        .b(stage0_col123[4]),
        .c_in(stage0_col123[5]),
        .s(fa_s0_c123_n962_s),
        .c_out(fa_s0_c123_n962_c)
    );

    fa fa_s0_c123_n963 (
        .a(stage0_col123[6]),
        .b(stage0_col123[7]),
        .c_in(stage0_col123[8]),
        .s(fa_s0_c123_n963_s),
        .c_out(fa_s0_c123_n963_c)
    );

    fa fa_s0_c123_n964 (
        .a(stage0_col123[9]),
        .b(stage0_col123[10]),
        .c_in(stage0_col123[11]),
        .s(fa_s0_c123_n964_s),
        .c_out(fa_s0_c123_n964_c)
    );

    fa fa_s0_c123_n965 (
        .a(stage0_col123[12]),
        .b(stage0_col123[13]),
        .c_in(stage0_col123[14]),
        .s(fa_s0_c123_n965_s),
        .c_out(fa_s0_c123_n965_c)
    );

    fa fa_s0_c123_n966 (
        .a(stage0_col123[15]),
        .b(stage0_col123[16]),
        .c_in(stage0_col123[17]),
        .s(fa_s0_c123_n966_s),
        .c_out(fa_s0_c123_n966_c)
    );

    fa fa_s0_c123_n967 (
        .a(stage0_col123[18]),
        .b(stage0_col123[19]),
        .c_in(stage0_col123[20]),
        .s(fa_s0_c123_n967_s),
        .c_out(fa_s0_c123_n967_c)
    );

    fa fa_s0_c123_n968 (
        .a(stage0_col123[21]),
        .b(stage0_col123[22]),
        .c_in(stage0_col123[23]),
        .s(fa_s0_c123_n968_s),
        .c_out(fa_s0_c123_n968_c)
    );

    fa fa_s0_c123_n969 (
        .a(stage0_col123[24]),
        .b(stage0_col123[25]),
        .c_in(stage0_col123[26]),
        .s(fa_s0_c123_n969_s),
        .c_out(fa_s0_c123_n969_c)
    );

    fa fa_s0_c123_n970 (
        .a(stage0_col123[27]),
        .b(stage0_col123[28]),
        .c_in(stage0_col123[29]),
        .s(fa_s0_c123_n970_s),
        .c_out(fa_s0_c123_n970_c)
    );

    fa fa_s0_c124_n971 (
        .a(stage0_col124[0]),
        .b(stage0_col124[1]),
        .c_in(stage0_col124[2]),
        .s(fa_s0_c124_n971_s),
        .c_out(fa_s0_c124_n971_c)
    );

    fa fa_s0_c124_n972 (
        .a(stage0_col124[3]),
        .b(stage0_col124[4]),
        .c_in(stage0_col124[5]),
        .s(fa_s0_c124_n972_s),
        .c_out(fa_s0_c124_n972_c)
    );

    fa fa_s0_c124_n973 (
        .a(stage0_col124[6]),
        .b(stage0_col124[7]),
        .c_in(stage0_col124[8]),
        .s(fa_s0_c124_n973_s),
        .c_out(fa_s0_c124_n973_c)
    );

    fa fa_s0_c124_n974 (
        .a(stage0_col124[9]),
        .b(stage0_col124[10]),
        .c_in(stage0_col124[11]),
        .s(fa_s0_c124_n974_s),
        .c_out(fa_s0_c124_n974_c)
    );

    fa fa_s0_c124_n975 (
        .a(stage0_col124[12]),
        .b(stage0_col124[13]),
        .c_in(stage0_col124[14]),
        .s(fa_s0_c124_n975_s),
        .c_out(fa_s0_c124_n975_c)
    );

    fa fa_s0_c124_n976 (
        .a(stage0_col124[15]),
        .b(stage0_col124[16]),
        .c_in(stage0_col124[17]),
        .s(fa_s0_c124_n976_s),
        .c_out(fa_s0_c124_n976_c)
    );

    fa fa_s0_c124_n977 (
        .a(stage0_col124[18]),
        .b(stage0_col124[19]),
        .c_in(stage0_col124[20]),
        .s(fa_s0_c124_n977_s),
        .c_out(fa_s0_c124_n977_c)
    );

    fa fa_s0_c124_n978 (
        .a(stage0_col124[21]),
        .b(stage0_col124[22]),
        .c_in(stage0_col124[23]),
        .s(fa_s0_c124_n978_s),
        .c_out(fa_s0_c124_n978_c)
    );

    fa fa_s0_c124_n979 (
        .a(stage0_col124[24]),
        .b(stage0_col124[25]),
        .c_in(stage0_col124[26]),
        .s(fa_s0_c124_n979_s),
        .c_out(fa_s0_c124_n979_c)
    );

    fa fa_s0_c124_n980 (
        .a(stage0_col124[27]),
        .b(stage0_col124[28]),
        .c_in(stage0_col124[29]),
        .s(fa_s0_c124_n980_s),
        .c_out(fa_s0_c124_n980_c)
    );

    fa fa_s0_c124_n981 (
        .a(stage0_col124[30]),
        .b(stage0_col124[31]),
        .c_in(stage0_col124[32]),
        .s(fa_s0_c124_n981_s),
        .c_out(fa_s0_c124_n981_c)
    );

    fa fa_s0_c125_n982 (
        .a(stage0_col125[0]),
        .b(stage0_col125[1]),
        .c_in(stage0_col125[2]),
        .s(fa_s0_c125_n982_s),
        .c_out(fa_s0_c125_n982_c)
    );

    fa fa_s0_c125_n983 (
        .a(stage0_col125[3]),
        .b(stage0_col125[4]),
        .c_in(stage0_col125[5]),
        .s(fa_s0_c125_n983_s),
        .c_out(fa_s0_c125_n983_c)
    );

    fa fa_s0_c125_n984 (
        .a(stage0_col125[6]),
        .b(stage0_col125[7]),
        .c_in(stage0_col125[8]),
        .s(fa_s0_c125_n984_s),
        .c_out(fa_s0_c125_n984_c)
    );

    fa fa_s0_c125_n985 (
        .a(stage0_col125[9]),
        .b(stage0_col125[10]),
        .c_in(stage0_col125[11]),
        .s(fa_s0_c125_n985_s),
        .c_out(fa_s0_c125_n985_c)
    );

    fa fa_s0_c125_n986 (
        .a(stage0_col125[12]),
        .b(stage0_col125[13]),
        .c_in(stage0_col125[14]),
        .s(fa_s0_c125_n986_s),
        .c_out(fa_s0_c125_n986_c)
    );

    fa fa_s0_c125_n987 (
        .a(stage0_col125[15]),
        .b(stage0_col125[16]),
        .c_in(stage0_col125[17]),
        .s(fa_s0_c125_n987_s),
        .c_out(fa_s0_c125_n987_c)
    );

    fa fa_s0_c125_n988 (
        .a(stage0_col125[18]),
        .b(stage0_col125[19]),
        .c_in(stage0_col125[20]),
        .s(fa_s0_c125_n988_s),
        .c_out(fa_s0_c125_n988_c)
    );

    fa fa_s0_c125_n989 (
        .a(stage0_col125[21]),
        .b(stage0_col125[22]),
        .c_in(stage0_col125[23]),
        .s(fa_s0_c125_n989_s),
        .c_out(fa_s0_c125_n989_c)
    );

    fa fa_s0_c125_n990 (
        .a(stage0_col125[24]),
        .b(stage0_col125[25]),
        .c_in(stage0_col125[26]),
        .s(fa_s0_c125_n990_s),
        .c_out(fa_s0_c125_n990_c)
    );

    fa fa_s0_c125_n991 (
        .a(stage0_col125[27]),
        .b(stage0_col125[28]),
        .c_in(stage0_col125[29]),
        .s(fa_s0_c125_n991_s),
        .c_out(fa_s0_c125_n991_c)
    );

    fa fa_s0_c126_n992 (
        .a(stage0_col126[0]),
        .b(stage0_col126[1]),
        .c_in(stage0_col126[2]),
        .s(fa_s0_c126_n992_s),
        .c_out(fa_s0_c126_n992_c)
    );

    fa fa_s0_c126_n993 (
        .a(stage0_col126[3]),
        .b(stage0_col126[4]),
        .c_in(stage0_col126[5]),
        .s(fa_s0_c126_n993_s),
        .c_out(fa_s0_c126_n993_c)
    );

    fa fa_s0_c126_n994 (
        .a(stage0_col126[6]),
        .b(stage0_col126[7]),
        .c_in(stage0_col126[8]),
        .s(fa_s0_c126_n994_s),
        .c_out(fa_s0_c126_n994_c)
    );

    fa fa_s0_c126_n995 (
        .a(stage0_col126[9]),
        .b(stage0_col126[10]),
        .c_in(stage0_col126[11]),
        .s(fa_s0_c126_n995_s),
        .c_out(fa_s0_c126_n995_c)
    );

    fa fa_s0_c126_n996 (
        .a(stage0_col126[12]),
        .b(stage0_col126[13]),
        .c_in(stage0_col126[14]),
        .s(fa_s0_c126_n996_s),
        .c_out(fa_s0_c126_n996_c)
    );

    fa fa_s0_c126_n997 (
        .a(stage0_col126[15]),
        .b(stage0_col126[16]),
        .c_in(stage0_col126[17]),
        .s(fa_s0_c126_n997_s),
        .c_out(fa_s0_c126_n997_c)
    );

    fa fa_s0_c126_n998 (
        .a(stage0_col126[18]),
        .b(stage0_col126[19]),
        .c_in(stage0_col126[20]),
        .s(fa_s0_c126_n998_s),
        .c_out(fa_s0_c126_n998_c)
    );

    fa fa_s0_c126_n999 (
        .a(stage0_col126[21]),
        .b(stage0_col126[22]),
        .c_in(stage0_col126[23]),
        .s(fa_s0_c126_n999_s),
        .c_out(fa_s0_c126_n999_c)
    );

    fa fa_s0_c126_n1000 (
        .a(stage0_col126[24]),
        .b(stage0_col126[25]),
        .c_in(stage0_col126[26]),
        .s(fa_s0_c126_n1000_s),
        .c_out(fa_s0_c126_n1000_c)
    );

    fa fa_s0_c126_n1001 (
        .a(stage0_col126[27]),
        .b(stage0_col126[28]),
        .c_in(stage0_col126[29]),
        .s(fa_s0_c126_n1001_s),
        .c_out(fa_s0_c126_n1001_c)
    );

    fa fa_s0_c126_n1002 (
        .a(stage0_col126[30]),
        .b(stage0_col126[31]),
        .c_in(stage0_col126[32]),
        .s(fa_s0_c126_n1002_s),
        .c_out(fa_s0_c126_n1002_c)
    );

    ha ha_s0_c0_n0 (
        .a(stage0_col0[0]),
        .b(stage0_col0[1]),
        .s(ha_s0_c0_n0_s),
        .c_out(ha_s0_c0_n0_c)
    );

    // Map to Stage 1 columns
    generate
        if (PIPE) begin : gen_stage1_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage1_col0[0] <= 1'b0;
                    stage1_col1[0] <= 1'b0;
                    stage1_col1[1] <= 1'b0;
                    stage1_col2[0] <= 1'b0;
                    stage1_col3[0] <= 1'b0;
                    stage1_col3[1] <= 1'b0;
                    stage1_col3[2] <= 1'b0;
                    stage1_col4[0] <= 1'b0;
                    stage1_col4[1] <= 1'b0;
                    stage1_col5[0] <= 1'b0;
                    stage1_col5[1] <= 1'b0;
                    stage1_col6[0] <= 1'b0;
                    stage1_col6[1] <= 1'b0;
                    stage1_col6[2] <= 1'b0;
                    stage1_col6[3] <= 1'b0;
                    stage1_col7[0] <= 1'b0;
                    stage1_col7[1] <= 1'b0;
                    stage1_col7[2] <= 1'b0;
                    stage1_col8[0] <= 1'b0;
                    stage1_col8[1] <= 1'b0;
                    stage1_col8[2] <= 1'b0;
                    stage1_col9[0] <= 1'b0;
                    stage1_col9[1] <= 1'b0;
                    stage1_col9[2] <= 1'b0;
                    stage1_col9[3] <= 1'b0;
                    stage1_col9[4] <= 1'b0;
                    stage1_col10[0] <= 1'b0;
                    stage1_col10[1] <= 1'b0;
                    stage1_col10[2] <= 1'b0;
                    stage1_col10[3] <= 1'b0;
                    stage1_col11[0] <= 1'b0;
                    stage1_col11[1] <= 1'b0;
                    stage1_col11[2] <= 1'b0;
                    stage1_col11[3] <= 1'b0;
                    stage1_col12[0] <= 1'b0;
                    stage1_col12[1] <= 1'b0;
                    stage1_col12[2] <= 1'b0;
                    stage1_col12[3] <= 1'b0;
                    stage1_col12[4] <= 1'b0;
                    stage1_col12[5] <= 1'b0;
                    stage1_col13[0] <= 1'b0;
                    stage1_col13[1] <= 1'b0;
                    stage1_col13[2] <= 1'b0;
                    stage1_col13[3] <= 1'b0;
                    stage1_col13[4] <= 1'b0;
                    stage1_col14[0] <= 1'b0;
                    stage1_col14[1] <= 1'b0;
                    stage1_col14[2] <= 1'b0;
                    stage1_col14[3] <= 1'b0;
                    stage1_col14[4] <= 1'b0;
                    stage1_col15[0] <= 1'b0;
                    stage1_col15[1] <= 1'b0;
                    stage1_col15[2] <= 1'b0;
                    stage1_col15[3] <= 1'b0;
                    stage1_col15[4] <= 1'b0;
                    stage1_col15[5] <= 1'b0;
                    stage1_col15[6] <= 1'b0;
                    stage1_col16[0] <= 1'b0;
                    stage1_col16[1] <= 1'b0;
                    stage1_col16[2] <= 1'b0;
                    stage1_col16[3] <= 1'b0;
                    stage1_col16[4] <= 1'b0;
                    stage1_col16[5] <= 1'b0;
                    stage1_col17[0] <= 1'b0;
                    stage1_col17[1] <= 1'b0;
                    stage1_col17[2] <= 1'b0;
                    stage1_col17[3] <= 1'b0;
                    stage1_col17[4] <= 1'b0;
                    stage1_col17[5] <= 1'b0;
                    stage1_col18[0] <= 1'b0;
                    stage1_col18[1] <= 1'b0;
                    stage1_col18[2] <= 1'b0;
                    stage1_col18[3] <= 1'b0;
                    stage1_col18[4] <= 1'b0;
                    stage1_col18[5] <= 1'b0;
                    stage1_col18[6] <= 1'b0;
                    stage1_col18[7] <= 1'b0;
                    stage1_col19[0] <= 1'b0;
                    stage1_col19[1] <= 1'b0;
                    stage1_col19[2] <= 1'b0;
                    stage1_col19[3] <= 1'b0;
                    stage1_col19[4] <= 1'b0;
                    stage1_col19[5] <= 1'b0;
                    stage1_col19[6] <= 1'b0;
                    stage1_col20[0] <= 1'b0;
                    stage1_col20[1] <= 1'b0;
                    stage1_col20[2] <= 1'b0;
                    stage1_col20[3] <= 1'b0;
                    stage1_col20[4] <= 1'b0;
                    stage1_col20[5] <= 1'b0;
                    stage1_col20[6] <= 1'b0;
                    stage1_col21[0] <= 1'b0;
                    stage1_col21[1] <= 1'b0;
                    stage1_col21[2] <= 1'b0;
                    stage1_col21[3] <= 1'b0;
                    stage1_col21[4] <= 1'b0;
                    stage1_col21[5] <= 1'b0;
                    stage1_col21[6] <= 1'b0;
                    stage1_col21[7] <= 1'b0;
                    stage1_col21[8] <= 1'b0;
                    stage1_col22[0] <= 1'b0;
                    stage1_col22[1] <= 1'b0;
                    stage1_col22[2] <= 1'b0;
                    stage1_col22[3] <= 1'b0;
                    stage1_col22[4] <= 1'b0;
                    stage1_col22[5] <= 1'b0;
                    stage1_col22[6] <= 1'b0;
                    stage1_col22[7] <= 1'b0;
                    stage1_col23[0] <= 1'b0;
                    stage1_col23[1] <= 1'b0;
                    stage1_col23[2] <= 1'b0;
                    stage1_col23[3] <= 1'b0;
                    stage1_col23[4] <= 1'b0;
                    stage1_col23[5] <= 1'b0;
                    stage1_col23[6] <= 1'b0;
                    stage1_col23[7] <= 1'b0;
                    stage1_col24[0] <= 1'b0;
                    stage1_col24[1] <= 1'b0;
                    stage1_col24[2] <= 1'b0;
                    stage1_col24[3] <= 1'b0;
                    stage1_col24[4] <= 1'b0;
                    stage1_col24[5] <= 1'b0;
                    stage1_col24[6] <= 1'b0;
                    stage1_col24[7] <= 1'b0;
                    stage1_col24[8] <= 1'b0;
                    stage1_col24[9] <= 1'b0;
                    stage1_col25[0] <= 1'b0;
                    stage1_col25[1] <= 1'b0;
                    stage1_col25[2] <= 1'b0;
                    stage1_col25[3] <= 1'b0;
                    stage1_col25[4] <= 1'b0;
                    stage1_col25[5] <= 1'b0;
                    stage1_col25[6] <= 1'b0;
                    stage1_col25[7] <= 1'b0;
                    stage1_col25[8] <= 1'b0;
                    stage1_col26[0] <= 1'b0;
                    stage1_col26[1] <= 1'b0;
                    stage1_col26[2] <= 1'b0;
                    stage1_col26[3] <= 1'b0;
                    stage1_col26[4] <= 1'b0;
                    stage1_col26[5] <= 1'b0;
                    stage1_col26[6] <= 1'b0;
                    stage1_col26[7] <= 1'b0;
                    stage1_col26[8] <= 1'b0;
                    stage1_col27[0] <= 1'b0;
                    stage1_col27[1] <= 1'b0;
                    stage1_col27[2] <= 1'b0;
                    stage1_col27[3] <= 1'b0;
                    stage1_col27[4] <= 1'b0;
                    stage1_col27[5] <= 1'b0;
                    stage1_col27[6] <= 1'b0;
                    stage1_col27[7] <= 1'b0;
                    stage1_col27[8] <= 1'b0;
                    stage1_col27[9] <= 1'b0;
                    stage1_col27[10] <= 1'b0;
                    stage1_col28[0] <= 1'b0;
                    stage1_col28[1] <= 1'b0;
                    stage1_col28[2] <= 1'b0;
                    stage1_col28[3] <= 1'b0;
                    stage1_col28[4] <= 1'b0;
                    stage1_col28[5] <= 1'b0;
                    stage1_col28[6] <= 1'b0;
                    stage1_col28[7] <= 1'b0;
                    stage1_col28[8] <= 1'b0;
                    stage1_col28[9] <= 1'b0;
                    stage1_col29[0] <= 1'b0;
                    stage1_col29[1] <= 1'b0;
                    stage1_col29[2] <= 1'b0;
                    stage1_col29[3] <= 1'b0;
                    stage1_col29[4] <= 1'b0;
                    stage1_col29[5] <= 1'b0;
                    stage1_col29[6] <= 1'b0;
                    stage1_col29[7] <= 1'b0;
                    stage1_col29[8] <= 1'b0;
                    stage1_col29[9] <= 1'b0;
                    stage1_col30[0] <= 1'b0;
                    stage1_col30[1] <= 1'b0;
                    stage1_col30[2] <= 1'b0;
                    stage1_col30[3] <= 1'b0;
                    stage1_col30[4] <= 1'b0;
                    stage1_col30[5] <= 1'b0;
                    stage1_col30[6] <= 1'b0;
                    stage1_col30[7] <= 1'b0;
                    stage1_col30[8] <= 1'b0;
                    stage1_col30[9] <= 1'b0;
                    stage1_col30[10] <= 1'b0;
                    stage1_col30[11] <= 1'b0;
                    stage1_col31[0] <= 1'b0;
                    stage1_col31[1] <= 1'b0;
                    stage1_col31[2] <= 1'b0;
                    stage1_col31[3] <= 1'b0;
                    stage1_col31[4] <= 1'b0;
                    stage1_col31[5] <= 1'b0;
                    stage1_col31[6] <= 1'b0;
                    stage1_col31[7] <= 1'b0;
                    stage1_col31[8] <= 1'b0;
                    stage1_col31[9] <= 1'b0;
                    stage1_col31[10] <= 1'b0;
                    stage1_col32[0] <= 1'b0;
                    stage1_col32[1] <= 1'b0;
                    stage1_col32[2] <= 1'b0;
                    stage1_col32[3] <= 1'b0;
                    stage1_col32[4] <= 1'b0;
                    stage1_col32[5] <= 1'b0;
                    stage1_col32[6] <= 1'b0;
                    stage1_col32[7] <= 1'b0;
                    stage1_col32[8] <= 1'b0;
                    stage1_col32[9] <= 1'b0;
                    stage1_col32[10] <= 1'b0;
                    stage1_col33[0] <= 1'b0;
                    stage1_col33[1] <= 1'b0;
                    stage1_col33[2] <= 1'b0;
                    stage1_col33[3] <= 1'b0;
                    stage1_col33[4] <= 1'b0;
                    stage1_col33[5] <= 1'b0;
                    stage1_col33[6] <= 1'b0;
                    stage1_col33[7] <= 1'b0;
                    stage1_col33[8] <= 1'b0;
                    stage1_col33[9] <= 1'b0;
                    stage1_col33[10] <= 1'b0;
                    stage1_col33[11] <= 1'b0;
                    stage1_col33[12] <= 1'b0;
                    stage1_col34[0] <= 1'b0;
                    stage1_col34[1] <= 1'b0;
                    stage1_col34[2] <= 1'b0;
                    stage1_col34[3] <= 1'b0;
                    stage1_col34[4] <= 1'b0;
                    stage1_col34[5] <= 1'b0;
                    stage1_col34[6] <= 1'b0;
                    stage1_col34[7] <= 1'b0;
                    stage1_col34[8] <= 1'b0;
                    stage1_col34[9] <= 1'b0;
                    stage1_col34[10] <= 1'b0;
                    stage1_col34[11] <= 1'b0;
                    stage1_col35[0] <= 1'b0;
                    stage1_col35[1] <= 1'b0;
                    stage1_col35[2] <= 1'b0;
                    stage1_col35[3] <= 1'b0;
                    stage1_col35[4] <= 1'b0;
                    stage1_col35[5] <= 1'b0;
                    stage1_col35[6] <= 1'b0;
                    stage1_col35[7] <= 1'b0;
                    stage1_col35[8] <= 1'b0;
                    stage1_col35[9] <= 1'b0;
                    stage1_col35[10] <= 1'b0;
                    stage1_col35[11] <= 1'b0;
                    stage1_col36[0] <= 1'b0;
                    stage1_col36[1] <= 1'b0;
                    stage1_col36[2] <= 1'b0;
                    stage1_col36[3] <= 1'b0;
                    stage1_col36[4] <= 1'b0;
                    stage1_col36[5] <= 1'b0;
                    stage1_col36[6] <= 1'b0;
                    stage1_col36[7] <= 1'b0;
                    stage1_col36[8] <= 1'b0;
                    stage1_col36[9] <= 1'b0;
                    stage1_col36[10] <= 1'b0;
                    stage1_col36[11] <= 1'b0;
                    stage1_col36[12] <= 1'b0;
                    stage1_col36[13] <= 1'b0;
                    stage1_col37[0] <= 1'b0;
                    stage1_col37[1] <= 1'b0;
                    stage1_col37[2] <= 1'b0;
                    stage1_col37[3] <= 1'b0;
                    stage1_col37[4] <= 1'b0;
                    stage1_col37[5] <= 1'b0;
                    stage1_col37[6] <= 1'b0;
                    stage1_col37[7] <= 1'b0;
                    stage1_col37[8] <= 1'b0;
                    stage1_col37[9] <= 1'b0;
                    stage1_col37[10] <= 1'b0;
                    stage1_col37[11] <= 1'b0;
                    stage1_col37[12] <= 1'b0;
                    stage1_col38[0] <= 1'b0;
                    stage1_col38[1] <= 1'b0;
                    stage1_col38[2] <= 1'b0;
                    stage1_col38[3] <= 1'b0;
                    stage1_col38[4] <= 1'b0;
                    stage1_col38[5] <= 1'b0;
                    stage1_col38[6] <= 1'b0;
                    stage1_col38[7] <= 1'b0;
                    stage1_col38[8] <= 1'b0;
                    stage1_col38[9] <= 1'b0;
                    stage1_col38[10] <= 1'b0;
                    stage1_col38[11] <= 1'b0;
                    stage1_col38[12] <= 1'b0;
                    stage1_col39[0] <= 1'b0;
                    stage1_col39[1] <= 1'b0;
                    stage1_col39[2] <= 1'b0;
                    stage1_col39[3] <= 1'b0;
                    stage1_col39[4] <= 1'b0;
                    stage1_col39[5] <= 1'b0;
                    stage1_col39[6] <= 1'b0;
                    stage1_col39[7] <= 1'b0;
                    stage1_col39[8] <= 1'b0;
                    stage1_col39[9] <= 1'b0;
                    stage1_col39[10] <= 1'b0;
                    stage1_col39[11] <= 1'b0;
                    stage1_col39[12] <= 1'b0;
                    stage1_col39[13] <= 1'b0;
                    stage1_col39[14] <= 1'b0;
                    stage1_col40[0] <= 1'b0;
                    stage1_col40[1] <= 1'b0;
                    stage1_col40[2] <= 1'b0;
                    stage1_col40[3] <= 1'b0;
                    stage1_col40[4] <= 1'b0;
                    stage1_col40[5] <= 1'b0;
                    stage1_col40[6] <= 1'b0;
                    stage1_col40[7] <= 1'b0;
                    stage1_col40[8] <= 1'b0;
                    stage1_col40[9] <= 1'b0;
                    stage1_col40[10] <= 1'b0;
                    stage1_col40[11] <= 1'b0;
                    stage1_col40[12] <= 1'b0;
                    stage1_col40[13] <= 1'b0;
                    stage1_col41[0] <= 1'b0;
                    stage1_col41[1] <= 1'b0;
                    stage1_col41[2] <= 1'b0;
                    stage1_col41[3] <= 1'b0;
                    stage1_col41[4] <= 1'b0;
                    stage1_col41[5] <= 1'b0;
                    stage1_col41[6] <= 1'b0;
                    stage1_col41[7] <= 1'b0;
                    stage1_col41[8] <= 1'b0;
                    stage1_col41[9] <= 1'b0;
                    stage1_col41[10] <= 1'b0;
                    stage1_col41[11] <= 1'b0;
                    stage1_col41[12] <= 1'b0;
                    stage1_col41[13] <= 1'b0;
                    stage1_col42[0] <= 1'b0;
                    stage1_col42[1] <= 1'b0;
                    stage1_col42[2] <= 1'b0;
                    stage1_col42[3] <= 1'b0;
                    stage1_col42[4] <= 1'b0;
                    stage1_col42[5] <= 1'b0;
                    stage1_col42[6] <= 1'b0;
                    stage1_col42[7] <= 1'b0;
                    stage1_col42[8] <= 1'b0;
                    stage1_col42[9] <= 1'b0;
                    stage1_col42[10] <= 1'b0;
                    stage1_col42[11] <= 1'b0;
                    stage1_col42[12] <= 1'b0;
                    stage1_col42[13] <= 1'b0;
                    stage1_col42[14] <= 1'b0;
                    stage1_col42[15] <= 1'b0;
                    stage1_col43[0] <= 1'b0;
                    stage1_col43[1] <= 1'b0;
                    stage1_col43[2] <= 1'b0;
                    stage1_col43[3] <= 1'b0;
                    stage1_col43[4] <= 1'b0;
                    stage1_col43[5] <= 1'b0;
                    stage1_col43[6] <= 1'b0;
                    stage1_col43[7] <= 1'b0;
                    stage1_col43[8] <= 1'b0;
                    stage1_col43[9] <= 1'b0;
                    stage1_col43[10] <= 1'b0;
                    stage1_col43[11] <= 1'b0;
                    stage1_col43[12] <= 1'b0;
                    stage1_col43[13] <= 1'b0;
                    stage1_col43[14] <= 1'b0;
                    stage1_col44[0] <= 1'b0;
                    stage1_col44[1] <= 1'b0;
                    stage1_col44[2] <= 1'b0;
                    stage1_col44[3] <= 1'b0;
                    stage1_col44[4] <= 1'b0;
                    stage1_col44[5] <= 1'b0;
                    stage1_col44[6] <= 1'b0;
                    stage1_col44[7] <= 1'b0;
                    stage1_col44[8] <= 1'b0;
                    stage1_col44[9] <= 1'b0;
                    stage1_col44[10] <= 1'b0;
                    stage1_col44[11] <= 1'b0;
                    stage1_col44[12] <= 1'b0;
                    stage1_col44[13] <= 1'b0;
                    stage1_col44[14] <= 1'b0;
                    stage1_col45[0] <= 1'b0;
                    stage1_col45[1] <= 1'b0;
                    stage1_col45[2] <= 1'b0;
                    stage1_col45[3] <= 1'b0;
                    stage1_col45[4] <= 1'b0;
                    stage1_col45[5] <= 1'b0;
                    stage1_col45[6] <= 1'b0;
                    stage1_col45[7] <= 1'b0;
                    stage1_col45[8] <= 1'b0;
                    stage1_col45[9] <= 1'b0;
                    stage1_col45[10] <= 1'b0;
                    stage1_col45[11] <= 1'b0;
                    stage1_col45[12] <= 1'b0;
                    stage1_col45[13] <= 1'b0;
                    stage1_col45[14] <= 1'b0;
                    stage1_col45[15] <= 1'b0;
                    stage1_col45[16] <= 1'b0;
                    stage1_col46[0] <= 1'b0;
                    stage1_col46[1] <= 1'b0;
                    stage1_col46[2] <= 1'b0;
                    stage1_col46[3] <= 1'b0;
                    stage1_col46[4] <= 1'b0;
                    stage1_col46[5] <= 1'b0;
                    stage1_col46[6] <= 1'b0;
                    stage1_col46[7] <= 1'b0;
                    stage1_col46[8] <= 1'b0;
                    stage1_col46[9] <= 1'b0;
                    stage1_col46[10] <= 1'b0;
                    stage1_col46[11] <= 1'b0;
                    stage1_col46[12] <= 1'b0;
                    stage1_col46[13] <= 1'b0;
                    stage1_col46[14] <= 1'b0;
                    stage1_col46[15] <= 1'b0;
                    stage1_col47[0] <= 1'b0;
                    stage1_col47[1] <= 1'b0;
                    stage1_col47[2] <= 1'b0;
                    stage1_col47[3] <= 1'b0;
                    stage1_col47[4] <= 1'b0;
                    stage1_col47[5] <= 1'b0;
                    stage1_col47[6] <= 1'b0;
                    stage1_col47[7] <= 1'b0;
                    stage1_col47[8] <= 1'b0;
                    stage1_col47[9] <= 1'b0;
                    stage1_col47[10] <= 1'b0;
                    stage1_col47[11] <= 1'b0;
                    stage1_col47[12] <= 1'b0;
                    stage1_col47[13] <= 1'b0;
                    stage1_col47[14] <= 1'b0;
                    stage1_col47[15] <= 1'b0;
                    stage1_col48[0] <= 1'b0;
                    stage1_col48[1] <= 1'b0;
                    stage1_col48[2] <= 1'b0;
                    stage1_col48[3] <= 1'b0;
                    stage1_col48[4] <= 1'b0;
                    stage1_col48[5] <= 1'b0;
                    stage1_col48[6] <= 1'b0;
                    stage1_col48[7] <= 1'b0;
                    stage1_col48[8] <= 1'b0;
                    stage1_col48[9] <= 1'b0;
                    stage1_col48[10] <= 1'b0;
                    stage1_col48[11] <= 1'b0;
                    stage1_col48[12] <= 1'b0;
                    stage1_col48[13] <= 1'b0;
                    stage1_col48[14] <= 1'b0;
                    stage1_col48[15] <= 1'b0;
                    stage1_col48[16] <= 1'b0;
                    stage1_col48[17] <= 1'b0;
                    stage1_col49[0] <= 1'b0;
                    stage1_col49[1] <= 1'b0;
                    stage1_col49[2] <= 1'b0;
                    stage1_col49[3] <= 1'b0;
                    stage1_col49[4] <= 1'b0;
                    stage1_col49[5] <= 1'b0;
                    stage1_col49[6] <= 1'b0;
                    stage1_col49[7] <= 1'b0;
                    stage1_col49[8] <= 1'b0;
                    stage1_col49[9] <= 1'b0;
                    stage1_col49[10] <= 1'b0;
                    stage1_col49[11] <= 1'b0;
                    stage1_col49[12] <= 1'b0;
                    stage1_col49[13] <= 1'b0;
                    stage1_col49[14] <= 1'b0;
                    stage1_col49[15] <= 1'b0;
                    stage1_col49[16] <= 1'b0;
                    stage1_col50[0] <= 1'b0;
                    stage1_col50[1] <= 1'b0;
                    stage1_col50[2] <= 1'b0;
                    stage1_col50[3] <= 1'b0;
                    stage1_col50[4] <= 1'b0;
                    stage1_col50[5] <= 1'b0;
                    stage1_col50[6] <= 1'b0;
                    stage1_col50[7] <= 1'b0;
                    stage1_col50[8] <= 1'b0;
                    stage1_col50[9] <= 1'b0;
                    stage1_col50[10] <= 1'b0;
                    stage1_col50[11] <= 1'b0;
                    stage1_col50[12] <= 1'b0;
                    stage1_col50[13] <= 1'b0;
                    stage1_col50[14] <= 1'b0;
                    stage1_col50[15] <= 1'b0;
                    stage1_col50[16] <= 1'b0;
                    stage1_col51[0] <= 1'b0;
                    stage1_col51[1] <= 1'b0;
                    stage1_col51[2] <= 1'b0;
                    stage1_col51[3] <= 1'b0;
                    stage1_col51[4] <= 1'b0;
                    stage1_col51[5] <= 1'b0;
                    stage1_col51[6] <= 1'b0;
                    stage1_col51[7] <= 1'b0;
                    stage1_col51[8] <= 1'b0;
                    stage1_col51[9] <= 1'b0;
                    stage1_col51[10] <= 1'b0;
                    stage1_col51[11] <= 1'b0;
                    stage1_col51[12] <= 1'b0;
                    stage1_col51[13] <= 1'b0;
                    stage1_col51[14] <= 1'b0;
                    stage1_col51[15] <= 1'b0;
                    stage1_col51[16] <= 1'b0;
                    stage1_col51[17] <= 1'b0;
                    stage1_col51[18] <= 1'b0;
                    stage1_col52[0] <= 1'b0;
                    stage1_col52[1] <= 1'b0;
                    stage1_col52[2] <= 1'b0;
                    stage1_col52[3] <= 1'b0;
                    stage1_col52[4] <= 1'b0;
                    stage1_col52[5] <= 1'b0;
                    stage1_col52[6] <= 1'b0;
                    stage1_col52[7] <= 1'b0;
                    stage1_col52[8] <= 1'b0;
                    stage1_col52[9] <= 1'b0;
                    stage1_col52[10] <= 1'b0;
                    stage1_col52[11] <= 1'b0;
                    stage1_col52[12] <= 1'b0;
                    stage1_col52[13] <= 1'b0;
                    stage1_col52[14] <= 1'b0;
                    stage1_col52[15] <= 1'b0;
                    stage1_col52[16] <= 1'b0;
                    stage1_col52[17] <= 1'b0;
                    stage1_col53[0] <= 1'b0;
                    stage1_col53[1] <= 1'b0;
                    stage1_col53[2] <= 1'b0;
                    stage1_col53[3] <= 1'b0;
                    stage1_col53[4] <= 1'b0;
                    stage1_col53[5] <= 1'b0;
                    stage1_col53[6] <= 1'b0;
                    stage1_col53[7] <= 1'b0;
                    stage1_col53[8] <= 1'b0;
                    stage1_col53[9] <= 1'b0;
                    stage1_col53[10] <= 1'b0;
                    stage1_col53[11] <= 1'b0;
                    stage1_col53[12] <= 1'b0;
                    stage1_col53[13] <= 1'b0;
                    stage1_col53[14] <= 1'b0;
                    stage1_col53[15] <= 1'b0;
                    stage1_col53[16] <= 1'b0;
                    stage1_col53[17] <= 1'b0;
                    stage1_col54[0] <= 1'b0;
                    stage1_col54[1] <= 1'b0;
                    stage1_col54[2] <= 1'b0;
                    stage1_col54[3] <= 1'b0;
                    stage1_col54[4] <= 1'b0;
                    stage1_col54[5] <= 1'b0;
                    stage1_col54[6] <= 1'b0;
                    stage1_col54[7] <= 1'b0;
                    stage1_col54[8] <= 1'b0;
                    stage1_col54[9] <= 1'b0;
                    stage1_col54[10] <= 1'b0;
                    stage1_col54[11] <= 1'b0;
                    stage1_col54[12] <= 1'b0;
                    stage1_col54[13] <= 1'b0;
                    stage1_col54[14] <= 1'b0;
                    stage1_col54[15] <= 1'b0;
                    stage1_col54[16] <= 1'b0;
                    stage1_col54[17] <= 1'b0;
                    stage1_col54[18] <= 1'b0;
                    stage1_col54[19] <= 1'b0;
                    stage1_col55[0] <= 1'b0;
                    stage1_col55[1] <= 1'b0;
                    stage1_col55[2] <= 1'b0;
                    stage1_col55[3] <= 1'b0;
                    stage1_col55[4] <= 1'b0;
                    stage1_col55[5] <= 1'b0;
                    stage1_col55[6] <= 1'b0;
                    stage1_col55[7] <= 1'b0;
                    stage1_col55[8] <= 1'b0;
                    stage1_col55[9] <= 1'b0;
                    stage1_col55[10] <= 1'b0;
                    stage1_col55[11] <= 1'b0;
                    stage1_col55[12] <= 1'b0;
                    stage1_col55[13] <= 1'b0;
                    stage1_col55[14] <= 1'b0;
                    stage1_col55[15] <= 1'b0;
                    stage1_col55[16] <= 1'b0;
                    stage1_col55[17] <= 1'b0;
                    stage1_col55[18] <= 1'b0;
                    stage1_col56[0] <= 1'b0;
                    stage1_col56[1] <= 1'b0;
                    stage1_col56[2] <= 1'b0;
                    stage1_col56[3] <= 1'b0;
                    stage1_col56[4] <= 1'b0;
                    stage1_col56[5] <= 1'b0;
                    stage1_col56[6] <= 1'b0;
                    stage1_col56[7] <= 1'b0;
                    stage1_col56[8] <= 1'b0;
                    stage1_col56[9] <= 1'b0;
                    stage1_col56[10] <= 1'b0;
                    stage1_col56[11] <= 1'b0;
                    stage1_col56[12] <= 1'b0;
                    stage1_col56[13] <= 1'b0;
                    stage1_col56[14] <= 1'b0;
                    stage1_col56[15] <= 1'b0;
                    stage1_col56[16] <= 1'b0;
                    stage1_col56[17] <= 1'b0;
                    stage1_col56[18] <= 1'b0;
                    stage1_col57[0] <= 1'b0;
                    stage1_col57[1] <= 1'b0;
                    stage1_col57[2] <= 1'b0;
                    stage1_col57[3] <= 1'b0;
                    stage1_col57[4] <= 1'b0;
                    stage1_col57[5] <= 1'b0;
                    stage1_col57[6] <= 1'b0;
                    stage1_col57[7] <= 1'b0;
                    stage1_col57[8] <= 1'b0;
                    stage1_col57[9] <= 1'b0;
                    stage1_col57[10] <= 1'b0;
                    stage1_col57[11] <= 1'b0;
                    stage1_col57[12] <= 1'b0;
                    stage1_col57[13] <= 1'b0;
                    stage1_col57[14] <= 1'b0;
                    stage1_col57[15] <= 1'b0;
                    stage1_col57[16] <= 1'b0;
                    stage1_col57[17] <= 1'b0;
                    stage1_col57[18] <= 1'b0;
                    stage1_col57[19] <= 1'b0;
                    stage1_col57[20] <= 1'b0;
                    stage1_col58[0] <= 1'b0;
                    stage1_col58[1] <= 1'b0;
                    stage1_col58[2] <= 1'b0;
                    stage1_col58[3] <= 1'b0;
                    stage1_col58[4] <= 1'b0;
                    stage1_col58[5] <= 1'b0;
                    stage1_col58[6] <= 1'b0;
                    stage1_col58[7] <= 1'b0;
                    stage1_col58[8] <= 1'b0;
                    stage1_col58[9] <= 1'b0;
                    stage1_col58[10] <= 1'b0;
                    stage1_col58[11] <= 1'b0;
                    stage1_col58[12] <= 1'b0;
                    stage1_col58[13] <= 1'b0;
                    stage1_col58[14] <= 1'b0;
                    stage1_col58[15] <= 1'b0;
                    stage1_col58[16] <= 1'b0;
                    stage1_col58[17] <= 1'b0;
                    stage1_col58[18] <= 1'b0;
                    stage1_col58[19] <= 1'b0;
                    stage1_col59[0] <= 1'b0;
                    stage1_col59[1] <= 1'b0;
                    stage1_col59[2] <= 1'b0;
                    stage1_col59[3] <= 1'b0;
                    stage1_col59[4] <= 1'b0;
                    stage1_col59[5] <= 1'b0;
                    stage1_col59[6] <= 1'b0;
                    stage1_col59[7] <= 1'b0;
                    stage1_col59[8] <= 1'b0;
                    stage1_col59[9] <= 1'b0;
                    stage1_col59[10] <= 1'b0;
                    stage1_col59[11] <= 1'b0;
                    stage1_col59[12] <= 1'b0;
                    stage1_col59[13] <= 1'b0;
                    stage1_col59[14] <= 1'b0;
                    stage1_col59[15] <= 1'b0;
                    stage1_col59[16] <= 1'b0;
                    stage1_col59[17] <= 1'b0;
                    stage1_col59[18] <= 1'b0;
                    stage1_col59[19] <= 1'b0;
                    stage1_col60[0] <= 1'b0;
                    stage1_col60[1] <= 1'b0;
                    stage1_col60[2] <= 1'b0;
                    stage1_col60[3] <= 1'b0;
                    stage1_col60[4] <= 1'b0;
                    stage1_col60[5] <= 1'b0;
                    stage1_col60[6] <= 1'b0;
                    stage1_col60[7] <= 1'b0;
                    stage1_col60[8] <= 1'b0;
                    stage1_col60[9] <= 1'b0;
                    stage1_col60[10] <= 1'b0;
                    stage1_col60[11] <= 1'b0;
                    stage1_col60[12] <= 1'b0;
                    stage1_col60[13] <= 1'b0;
                    stage1_col60[14] <= 1'b0;
                    stage1_col60[15] <= 1'b0;
                    stage1_col60[16] <= 1'b0;
                    stage1_col60[17] <= 1'b0;
                    stage1_col60[18] <= 1'b0;
                    stage1_col60[19] <= 1'b0;
                    stage1_col60[20] <= 1'b0;
                    stage1_col60[21] <= 1'b0;
                    stage1_col61[0] <= 1'b0;
                    stage1_col61[1] <= 1'b0;
                    stage1_col61[2] <= 1'b0;
                    stage1_col61[3] <= 1'b0;
                    stage1_col61[4] <= 1'b0;
                    stage1_col61[5] <= 1'b0;
                    stage1_col61[6] <= 1'b0;
                    stage1_col61[7] <= 1'b0;
                    stage1_col61[8] <= 1'b0;
                    stage1_col61[9] <= 1'b0;
                    stage1_col61[10] <= 1'b0;
                    stage1_col61[11] <= 1'b0;
                    stage1_col61[12] <= 1'b0;
                    stage1_col61[13] <= 1'b0;
                    stage1_col61[14] <= 1'b0;
                    stage1_col61[15] <= 1'b0;
                    stage1_col61[16] <= 1'b0;
                    stage1_col61[17] <= 1'b0;
                    stage1_col61[18] <= 1'b0;
                    stage1_col61[19] <= 1'b0;
                    stage1_col61[20] <= 1'b0;
                    stage1_col62[0] <= 1'b0;
                    stage1_col62[1] <= 1'b0;
                    stage1_col62[2] <= 1'b0;
                    stage1_col62[3] <= 1'b0;
                    stage1_col62[4] <= 1'b0;
                    stage1_col62[5] <= 1'b0;
                    stage1_col62[6] <= 1'b0;
                    stage1_col62[7] <= 1'b0;
                    stage1_col62[8] <= 1'b0;
                    stage1_col62[9] <= 1'b0;
                    stage1_col62[10] <= 1'b0;
                    stage1_col62[11] <= 1'b0;
                    stage1_col62[12] <= 1'b0;
                    stage1_col62[13] <= 1'b0;
                    stage1_col62[14] <= 1'b0;
                    stage1_col62[15] <= 1'b0;
                    stage1_col62[16] <= 1'b0;
                    stage1_col62[17] <= 1'b0;
                    stage1_col62[18] <= 1'b0;
                    stage1_col62[19] <= 1'b0;
                    stage1_col62[20] <= 1'b0;
                    stage1_col63[0] <= 1'b0;
                    stage1_col63[1] <= 1'b0;
                    stage1_col63[2] <= 1'b0;
                    stage1_col63[3] <= 1'b0;
                    stage1_col63[4] <= 1'b0;
                    stage1_col63[5] <= 1'b0;
                    stage1_col63[6] <= 1'b0;
                    stage1_col63[7] <= 1'b0;
                    stage1_col63[8] <= 1'b0;
                    stage1_col63[9] <= 1'b0;
                    stage1_col63[10] <= 1'b0;
                    stage1_col63[11] <= 1'b0;
                    stage1_col63[12] <= 1'b0;
                    stage1_col63[13] <= 1'b0;
                    stage1_col63[14] <= 1'b0;
                    stage1_col63[15] <= 1'b0;
                    stage1_col63[16] <= 1'b0;
                    stage1_col63[17] <= 1'b0;
                    stage1_col63[18] <= 1'b0;
                    stage1_col63[19] <= 1'b0;
                    stage1_col63[20] <= 1'b0;
                    stage1_col63[21] <= 1'b0;
                    stage1_col63[22] <= 1'b0;
                    stage1_col64[0] <= 1'b0;
                    stage1_col64[1] <= 1'b0;
                    stage1_col64[2] <= 1'b0;
                    stage1_col64[3] <= 1'b0;
                    stage1_col64[4] <= 1'b0;
                    stage1_col64[5] <= 1'b0;
                    stage1_col64[6] <= 1'b0;
                    stage1_col64[7] <= 1'b0;
                    stage1_col64[8] <= 1'b0;
                    stage1_col64[9] <= 1'b0;
                    stage1_col64[10] <= 1'b0;
                    stage1_col64[11] <= 1'b0;
                    stage1_col64[12] <= 1'b0;
                    stage1_col64[13] <= 1'b0;
                    stage1_col64[14] <= 1'b0;
                    stage1_col64[15] <= 1'b0;
                    stage1_col64[16] <= 1'b0;
                    stage1_col64[17] <= 1'b0;
                    stage1_col64[18] <= 1'b0;
                    stage1_col64[19] <= 1'b0;
                    stage1_col64[20] <= 1'b0;
                    stage1_col65[0] <= 1'b0;
                    stage1_col65[1] <= 1'b0;
                    stage1_col65[2] <= 1'b0;
                    stage1_col65[3] <= 1'b0;
                    stage1_col65[4] <= 1'b0;
                    stage1_col65[5] <= 1'b0;
                    stage1_col65[6] <= 1'b0;
                    stage1_col65[7] <= 1'b0;
                    stage1_col65[8] <= 1'b0;
                    stage1_col65[9] <= 1'b0;
                    stage1_col65[10] <= 1'b0;
                    stage1_col65[11] <= 1'b0;
                    stage1_col65[12] <= 1'b0;
                    stage1_col65[13] <= 1'b0;
                    stage1_col65[14] <= 1'b0;
                    stage1_col65[15] <= 1'b0;
                    stage1_col65[16] <= 1'b0;
                    stage1_col65[17] <= 1'b0;
                    stage1_col65[18] <= 1'b0;
                    stage1_col65[19] <= 1'b0;
                    stage1_col65[20] <= 1'b0;
                    stage1_col65[21] <= 1'b0;
                    stage1_col65[22] <= 1'b0;
                    stage1_col66[0] <= 1'b0;
                    stage1_col66[1] <= 1'b0;
                    stage1_col66[2] <= 1'b0;
                    stage1_col66[3] <= 1'b0;
                    stage1_col66[4] <= 1'b0;
                    stage1_col66[5] <= 1'b0;
                    stage1_col66[6] <= 1'b0;
                    stage1_col66[7] <= 1'b0;
                    stage1_col66[8] <= 1'b0;
                    stage1_col66[9] <= 1'b0;
                    stage1_col66[10] <= 1'b0;
                    stage1_col66[11] <= 1'b0;
                    stage1_col66[12] <= 1'b0;
                    stage1_col66[13] <= 1'b0;
                    stage1_col66[14] <= 1'b0;
                    stage1_col66[15] <= 1'b0;
                    stage1_col66[16] <= 1'b0;
                    stage1_col66[17] <= 1'b0;
                    stage1_col66[18] <= 1'b0;
                    stage1_col66[19] <= 1'b0;
                    stage1_col66[20] <= 1'b0;
                    stage1_col67[0] <= 1'b0;
                    stage1_col67[1] <= 1'b0;
                    stage1_col67[2] <= 1'b0;
                    stage1_col67[3] <= 1'b0;
                    stage1_col67[4] <= 1'b0;
                    stage1_col67[5] <= 1'b0;
                    stage1_col67[6] <= 1'b0;
                    stage1_col67[7] <= 1'b0;
                    stage1_col67[8] <= 1'b0;
                    stage1_col67[9] <= 1'b0;
                    stage1_col67[10] <= 1'b0;
                    stage1_col67[11] <= 1'b0;
                    stage1_col67[12] <= 1'b0;
                    stage1_col67[13] <= 1'b0;
                    stage1_col67[14] <= 1'b0;
                    stage1_col67[15] <= 1'b0;
                    stage1_col67[16] <= 1'b0;
                    stage1_col67[17] <= 1'b0;
                    stage1_col67[18] <= 1'b0;
                    stage1_col67[19] <= 1'b0;
                    stage1_col67[20] <= 1'b0;
                    stage1_col67[21] <= 1'b0;
                    stage1_col67[22] <= 1'b0;
                    stage1_col68[0] <= 1'b0;
                    stage1_col68[1] <= 1'b0;
                    stage1_col68[2] <= 1'b0;
                    stage1_col68[3] <= 1'b0;
                    stage1_col68[4] <= 1'b0;
                    stage1_col68[5] <= 1'b0;
                    stage1_col68[6] <= 1'b0;
                    stage1_col68[7] <= 1'b0;
                    stage1_col68[8] <= 1'b0;
                    stage1_col68[9] <= 1'b0;
                    stage1_col68[10] <= 1'b0;
                    stage1_col68[11] <= 1'b0;
                    stage1_col68[12] <= 1'b0;
                    stage1_col68[13] <= 1'b0;
                    stage1_col68[14] <= 1'b0;
                    stage1_col68[15] <= 1'b0;
                    stage1_col68[16] <= 1'b0;
                    stage1_col68[17] <= 1'b0;
                    stage1_col68[18] <= 1'b0;
                    stage1_col68[19] <= 1'b0;
                    stage1_col68[20] <= 1'b0;
                    stage1_col69[0] <= 1'b0;
                    stage1_col69[1] <= 1'b0;
                    stage1_col69[2] <= 1'b0;
                    stage1_col69[3] <= 1'b0;
                    stage1_col69[4] <= 1'b0;
                    stage1_col69[5] <= 1'b0;
                    stage1_col69[6] <= 1'b0;
                    stage1_col69[7] <= 1'b0;
                    stage1_col69[8] <= 1'b0;
                    stage1_col69[9] <= 1'b0;
                    stage1_col69[10] <= 1'b0;
                    stage1_col69[11] <= 1'b0;
                    stage1_col69[12] <= 1'b0;
                    stage1_col69[13] <= 1'b0;
                    stage1_col69[14] <= 1'b0;
                    stage1_col69[15] <= 1'b0;
                    stage1_col69[16] <= 1'b0;
                    stage1_col69[17] <= 1'b0;
                    stage1_col69[18] <= 1'b0;
                    stage1_col69[19] <= 1'b0;
                    stage1_col69[20] <= 1'b0;
                    stage1_col69[21] <= 1'b0;
                    stage1_col69[22] <= 1'b0;
                    stage1_col70[0] <= 1'b0;
                    stage1_col70[1] <= 1'b0;
                    stage1_col70[2] <= 1'b0;
                    stage1_col70[3] <= 1'b0;
                    stage1_col70[4] <= 1'b0;
                    stage1_col70[5] <= 1'b0;
                    stage1_col70[6] <= 1'b0;
                    stage1_col70[7] <= 1'b0;
                    stage1_col70[8] <= 1'b0;
                    stage1_col70[9] <= 1'b0;
                    stage1_col70[10] <= 1'b0;
                    stage1_col70[11] <= 1'b0;
                    stage1_col70[12] <= 1'b0;
                    stage1_col70[13] <= 1'b0;
                    stage1_col70[14] <= 1'b0;
                    stage1_col70[15] <= 1'b0;
                    stage1_col70[16] <= 1'b0;
                    stage1_col70[17] <= 1'b0;
                    stage1_col70[18] <= 1'b0;
                    stage1_col70[19] <= 1'b0;
                    stage1_col70[20] <= 1'b0;
                    stage1_col71[0] <= 1'b0;
                    stage1_col71[1] <= 1'b0;
                    stage1_col71[2] <= 1'b0;
                    stage1_col71[3] <= 1'b0;
                    stage1_col71[4] <= 1'b0;
                    stage1_col71[5] <= 1'b0;
                    stage1_col71[6] <= 1'b0;
                    stage1_col71[7] <= 1'b0;
                    stage1_col71[8] <= 1'b0;
                    stage1_col71[9] <= 1'b0;
                    stage1_col71[10] <= 1'b0;
                    stage1_col71[11] <= 1'b0;
                    stage1_col71[12] <= 1'b0;
                    stage1_col71[13] <= 1'b0;
                    stage1_col71[14] <= 1'b0;
                    stage1_col71[15] <= 1'b0;
                    stage1_col71[16] <= 1'b0;
                    stage1_col71[17] <= 1'b0;
                    stage1_col71[18] <= 1'b0;
                    stage1_col71[19] <= 1'b0;
                    stage1_col71[20] <= 1'b0;
                    stage1_col71[21] <= 1'b0;
                    stage1_col71[22] <= 1'b0;
                    stage1_col72[0] <= 1'b0;
                    stage1_col72[1] <= 1'b0;
                    stage1_col72[2] <= 1'b0;
                    stage1_col72[3] <= 1'b0;
                    stage1_col72[4] <= 1'b0;
                    stage1_col72[5] <= 1'b0;
                    stage1_col72[6] <= 1'b0;
                    stage1_col72[7] <= 1'b0;
                    stage1_col72[8] <= 1'b0;
                    stage1_col72[9] <= 1'b0;
                    stage1_col72[10] <= 1'b0;
                    stage1_col72[11] <= 1'b0;
                    stage1_col72[12] <= 1'b0;
                    stage1_col72[13] <= 1'b0;
                    stage1_col72[14] <= 1'b0;
                    stage1_col72[15] <= 1'b0;
                    stage1_col72[16] <= 1'b0;
                    stage1_col72[17] <= 1'b0;
                    stage1_col72[18] <= 1'b0;
                    stage1_col72[19] <= 1'b0;
                    stage1_col72[20] <= 1'b0;
                    stage1_col73[0] <= 1'b0;
                    stage1_col73[1] <= 1'b0;
                    stage1_col73[2] <= 1'b0;
                    stage1_col73[3] <= 1'b0;
                    stage1_col73[4] <= 1'b0;
                    stage1_col73[5] <= 1'b0;
                    stage1_col73[6] <= 1'b0;
                    stage1_col73[7] <= 1'b0;
                    stage1_col73[8] <= 1'b0;
                    stage1_col73[9] <= 1'b0;
                    stage1_col73[10] <= 1'b0;
                    stage1_col73[11] <= 1'b0;
                    stage1_col73[12] <= 1'b0;
                    stage1_col73[13] <= 1'b0;
                    stage1_col73[14] <= 1'b0;
                    stage1_col73[15] <= 1'b0;
                    stage1_col73[16] <= 1'b0;
                    stage1_col73[17] <= 1'b0;
                    stage1_col73[18] <= 1'b0;
                    stage1_col73[19] <= 1'b0;
                    stage1_col73[20] <= 1'b0;
                    stage1_col73[21] <= 1'b0;
                    stage1_col73[22] <= 1'b0;
                    stage1_col74[0] <= 1'b0;
                    stage1_col74[1] <= 1'b0;
                    stage1_col74[2] <= 1'b0;
                    stage1_col74[3] <= 1'b0;
                    stage1_col74[4] <= 1'b0;
                    stage1_col74[5] <= 1'b0;
                    stage1_col74[6] <= 1'b0;
                    stage1_col74[7] <= 1'b0;
                    stage1_col74[8] <= 1'b0;
                    stage1_col74[9] <= 1'b0;
                    stage1_col74[10] <= 1'b0;
                    stage1_col74[11] <= 1'b0;
                    stage1_col74[12] <= 1'b0;
                    stage1_col74[13] <= 1'b0;
                    stage1_col74[14] <= 1'b0;
                    stage1_col74[15] <= 1'b0;
                    stage1_col74[16] <= 1'b0;
                    stage1_col74[17] <= 1'b0;
                    stage1_col74[18] <= 1'b0;
                    stage1_col74[19] <= 1'b0;
                    stage1_col74[20] <= 1'b0;
                    stage1_col75[0] <= 1'b0;
                    stage1_col75[1] <= 1'b0;
                    stage1_col75[2] <= 1'b0;
                    stage1_col75[3] <= 1'b0;
                    stage1_col75[4] <= 1'b0;
                    stage1_col75[5] <= 1'b0;
                    stage1_col75[6] <= 1'b0;
                    stage1_col75[7] <= 1'b0;
                    stage1_col75[8] <= 1'b0;
                    stage1_col75[9] <= 1'b0;
                    stage1_col75[10] <= 1'b0;
                    stage1_col75[11] <= 1'b0;
                    stage1_col75[12] <= 1'b0;
                    stage1_col75[13] <= 1'b0;
                    stage1_col75[14] <= 1'b0;
                    stage1_col75[15] <= 1'b0;
                    stage1_col75[16] <= 1'b0;
                    stage1_col75[17] <= 1'b0;
                    stage1_col75[18] <= 1'b0;
                    stage1_col75[19] <= 1'b0;
                    stage1_col75[20] <= 1'b0;
                    stage1_col75[21] <= 1'b0;
                    stage1_col75[22] <= 1'b0;
                    stage1_col76[0] <= 1'b0;
                    stage1_col76[1] <= 1'b0;
                    stage1_col76[2] <= 1'b0;
                    stage1_col76[3] <= 1'b0;
                    stage1_col76[4] <= 1'b0;
                    stage1_col76[5] <= 1'b0;
                    stage1_col76[6] <= 1'b0;
                    stage1_col76[7] <= 1'b0;
                    stage1_col76[8] <= 1'b0;
                    stage1_col76[9] <= 1'b0;
                    stage1_col76[10] <= 1'b0;
                    stage1_col76[11] <= 1'b0;
                    stage1_col76[12] <= 1'b0;
                    stage1_col76[13] <= 1'b0;
                    stage1_col76[14] <= 1'b0;
                    stage1_col76[15] <= 1'b0;
                    stage1_col76[16] <= 1'b0;
                    stage1_col76[17] <= 1'b0;
                    stage1_col76[18] <= 1'b0;
                    stage1_col76[19] <= 1'b0;
                    stage1_col76[20] <= 1'b0;
                    stage1_col77[0] <= 1'b0;
                    stage1_col77[1] <= 1'b0;
                    stage1_col77[2] <= 1'b0;
                    stage1_col77[3] <= 1'b0;
                    stage1_col77[4] <= 1'b0;
                    stage1_col77[5] <= 1'b0;
                    stage1_col77[6] <= 1'b0;
                    stage1_col77[7] <= 1'b0;
                    stage1_col77[8] <= 1'b0;
                    stage1_col77[9] <= 1'b0;
                    stage1_col77[10] <= 1'b0;
                    stage1_col77[11] <= 1'b0;
                    stage1_col77[12] <= 1'b0;
                    stage1_col77[13] <= 1'b0;
                    stage1_col77[14] <= 1'b0;
                    stage1_col77[15] <= 1'b0;
                    stage1_col77[16] <= 1'b0;
                    stage1_col77[17] <= 1'b0;
                    stage1_col77[18] <= 1'b0;
                    stage1_col77[19] <= 1'b0;
                    stage1_col77[20] <= 1'b0;
                    stage1_col77[21] <= 1'b0;
                    stage1_col77[22] <= 1'b0;
                    stage1_col78[0] <= 1'b0;
                    stage1_col78[1] <= 1'b0;
                    stage1_col78[2] <= 1'b0;
                    stage1_col78[3] <= 1'b0;
                    stage1_col78[4] <= 1'b0;
                    stage1_col78[5] <= 1'b0;
                    stage1_col78[6] <= 1'b0;
                    stage1_col78[7] <= 1'b0;
                    stage1_col78[8] <= 1'b0;
                    stage1_col78[9] <= 1'b0;
                    stage1_col78[10] <= 1'b0;
                    stage1_col78[11] <= 1'b0;
                    stage1_col78[12] <= 1'b0;
                    stage1_col78[13] <= 1'b0;
                    stage1_col78[14] <= 1'b0;
                    stage1_col78[15] <= 1'b0;
                    stage1_col78[16] <= 1'b0;
                    stage1_col78[17] <= 1'b0;
                    stage1_col78[18] <= 1'b0;
                    stage1_col78[19] <= 1'b0;
                    stage1_col78[20] <= 1'b0;
                    stage1_col79[0] <= 1'b0;
                    stage1_col79[1] <= 1'b0;
                    stage1_col79[2] <= 1'b0;
                    stage1_col79[3] <= 1'b0;
                    stage1_col79[4] <= 1'b0;
                    stage1_col79[5] <= 1'b0;
                    stage1_col79[6] <= 1'b0;
                    stage1_col79[7] <= 1'b0;
                    stage1_col79[8] <= 1'b0;
                    stage1_col79[9] <= 1'b0;
                    stage1_col79[10] <= 1'b0;
                    stage1_col79[11] <= 1'b0;
                    stage1_col79[12] <= 1'b0;
                    stage1_col79[13] <= 1'b0;
                    stage1_col79[14] <= 1'b0;
                    stage1_col79[15] <= 1'b0;
                    stage1_col79[16] <= 1'b0;
                    stage1_col79[17] <= 1'b0;
                    stage1_col79[18] <= 1'b0;
                    stage1_col79[19] <= 1'b0;
                    stage1_col79[20] <= 1'b0;
                    stage1_col79[21] <= 1'b0;
                    stage1_col79[22] <= 1'b0;
                    stage1_col80[0] <= 1'b0;
                    stage1_col80[1] <= 1'b0;
                    stage1_col80[2] <= 1'b0;
                    stage1_col80[3] <= 1'b0;
                    stage1_col80[4] <= 1'b0;
                    stage1_col80[5] <= 1'b0;
                    stage1_col80[6] <= 1'b0;
                    stage1_col80[7] <= 1'b0;
                    stage1_col80[8] <= 1'b0;
                    stage1_col80[9] <= 1'b0;
                    stage1_col80[10] <= 1'b0;
                    stage1_col80[11] <= 1'b0;
                    stage1_col80[12] <= 1'b0;
                    stage1_col80[13] <= 1'b0;
                    stage1_col80[14] <= 1'b0;
                    stage1_col80[15] <= 1'b0;
                    stage1_col80[16] <= 1'b0;
                    stage1_col80[17] <= 1'b0;
                    stage1_col80[18] <= 1'b0;
                    stage1_col80[19] <= 1'b0;
                    stage1_col80[20] <= 1'b0;
                    stage1_col81[0] <= 1'b0;
                    stage1_col81[1] <= 1'b0;
                    stage1_col81[2] <= 1'b0;
                    stage1_col81[3] <= 1'b0;
                    stage1_col81[4] <= 1'b0;
                    stage1_col81[5] <= 1'b0;
                    stage1_col81[6] <= 1'b0;
                    stage1_col81[7] <= 1'b0;
                    stage1_col81[8] <= 1'b0;
                    stage1_col81[9] <= 1'b0;
                    stage1_col81[10] <= 1'b0;
                    stage1_col81[11] <= 1'b0;
                    stage1_col81[12] <= 1'b0;
                    stage1_col81[13] <= 1'b0;
                    stage1_col81[14] <= 1'b0;
                    stage1_col81[15] <= 1'b0;
                    stage1_col81[16] <= 1'b0;
                    stage1_col81[17] <= 1'b0;
                    stage1_col81[18] <= 1'b0;
                    stage1_col81[19] <= 1'b0;
                    stage1_col81[20] <= 1'b0;
                    stage1_col81[21] <= 1'b0;
                    stage1_col81[22] <= 1'b0;
                    stage1_col82[0] <= 1'b0;
                    stage1_col82[1] <= 1'b0;
                    stage1_col82[2] <= 1'b0;
                    stage1_col82[3] <= 1'b0;
                    stage1_col82[4] <= 1'b0;
                    stage1_col82[5] <= 1'b0;
                    stage1_col82[6] <= 1'b0;
                    stage1_col82[7] <= 1'b0;
                    stage1_col82[8] <= 1'b0;
                    stage1_col82[9] <= 1'b0;
                    stage1_col82[10] <= 1'b0;
                    stage1_col82[11] <= 1'b0;
                    stage1_col82[12] <= 1'b0;
                    stage1_col82[13] <= 1'b0;
                    stage1_col82[14] <= 1'b0;
                    stage1_col82[15] <= 1'b0;
                    stage1_col82[16] <= 1'b0;
                    stage1_col82[17] <= 1'b0;
                    stage1_col82[18] <= 1'b0;
                    stage1_col82[19] <= 1'b0;
                    stage1_col82[20] <= 1'b0;
                    stage1_col83[0] <= 1'b0;
                    stage1_col83[1] <= 1'b0;
                    stage1_col83[2] <= 1'b0;
                    stage1_col83[3] <= 1'b0;
                    stage1_col83[4] <= 1'b0;
                    stage1_col83[5] <= 1'b0;
                    stage1_col83[6] <= 1'b0;
                    stage1_col83[7] <= 1'b0;
                    stage1_col83[8] <= 1'b0;
                    stage1_col83[9] <= 1'b0;
                    stage1_col83[10] <= 1'b0;
                    stage1_col83[11] <= 1'b0;
                    stage1_col83[12] <= 1'b0;
                    stage1_col83[13] <= 1'b0;
                    stage1_col83[14] <= 1'b0;
                    stage1_col83[15] <= 1'b0;
                    stage1_col83[16] <= 1'b0;
                    stage1_col83[17] <= 1'b0;
                    stage1_col83[18] <= 1'b0;
                    stage1_col83[19] <= 1'b0;
                    stage1_col83[20] <= 1'b0;
                    stage1_col83[21] <= 1'b0;
                    stage1_col83[22] <= 1'b0;
                    stage1_col84[0] <= 1'b0;
                    stage1_col84[1] <= 1'b0;
                    stage1_col84[2] <= 1'b0;
                    stage1_col84[3] <= 1'b0;
                    stage1_col84[4] <= 1'b0;
                    stage1_col84[5] <= 1'b0;
                    stage1_col84[6] <= 1'b0;
                    stage1_col84[7] <= 1'b0;
                    stage1_col84[8] <= 1'b0;
                    stage1_col84[9] <= 1'b0;
                    stage1_col84[10] <= 1'b0;
                    stage1_col84[11] <= 1'b0;
                    stage1_col84[12] <= 1'b0;
                    stage1_col84[13] <= 1'b0;
                    stage1_col84[14] <= 1'b0;
                    stage1_col84[15] <= 1'b0;
                    stage1_col84[16] <= 1'b0;
                    stage1_col84[17] <= 1'b0;
                    stage1_col84[18] <= 1'b0;
                    stage1_col84[19] <= 1'b0;
                    stage1_col84[20] <= 1'b0;
                    stage1_col85[0] <= 1'b0;
                    stage1_col85[1] <= 1'b0;
                    stage1_col85[2] <= 1'b0;
                    stage1_col85[3] <= 1'b0;
                    stage1_col85[4] <= 1'b0;
                    stage1_col85[5] <= 1'b0;
                    stage1_col85[6] <= 1'b0;
                    stage1_col85[7] <= 1'b0;
                    stage1_col85[8] <= 1'b0;
                    stage1_col85[9] <= 1'b0;
                    stage1_col85[10] <= 1'b0;
                    stage1_col85[11] <= 1'b0;
                    stage1_col85[12] <= 1'b0;
                    stage1_col85[13] <= 1'b0;
                    stage1_col85[14] <= 1'b0;
                    stage1_col85[15] <= 1'b0;
                    stage1_col85[16] <= 1'b0;
                    stage1_col85[17] <= 1'b0;
                    stage1_col85[18] <= 1'b0;
                    stage1_col85[19] <= 1'b0;
                    stage1_col85[20] <= 1'b0;
                    stage1_col85[21] <= 1'b0;
                    stage1_col85[22] <= 1'b0;
                    stage1_col86[0] <= 1'b0;
                    stage1_col86[1] <= 1'b0;
                    stage1_col86[2] <= 1'b0;
                    stage1_col86[3] <= 1'b0;
                    stage1_col86[4] <= 1'b0;
                    stage1_col86[5] <= 1'b0;
                    stage1_col86[6] <= 1'b0;
                    stage1_col86[7] <= 1'b0;
                    stage1_col86[8] <= 1'b0;
                    stage1_col86[9] <= 1'b0;
                    stage1_col86[10] <= 1'b0;
                    stage1_col86[11] <= 1'b0;
                    stage1_col86[12] <= 1'b0;
                    stage1_col86[13] <= 1'b0;
                    stage1_col86[14] <= 1'b0;
                    stage1_col86[15] <= 1'b0;
                    stage1_col86[16] <= 1'b0;
                    stage1_col86[17] <= 1'b0;
                    stage1_col86[18] <= 1'b0;
                    stage1_col86[19] <= 1'b0;
                    stage1_col86[20] <= 1'b0;
                    stage1_col87[0] <= 1'b0;
                    stage1_col87[1] <= 1'b0;
                    stage1_col87[2] <= 1'b0;
                    stage1_col87[3] <= 1'b0;
                    stage1_col87[4] <= 1'b0;
                    stage1_col87[5] <= 1'b0;
                    stage1_col87[6] <= 1'b0;
                    stage1_col87[7] <= 1'b0;
                    stage1_col87[8] <= 1'b0;
                    stage1_col87[9] <= 1'b0;
                    stage1_col87[10] <= 1'b0;
                    stage1_col87[11] <= 1'b0;
                    stage1_col87[12] <= 1'b0;
                    stage1_col87[13] <= 1'b0;
                    stage1_col87[14] <= 1'b0;
                    stage1_col87[15] <= 1'b0;
                    stage1_col87[16] <= 1'b0;
                    stage1_col87[17] <= 1'b0;
                    stage1_col87[18] <= 1'b0;
                    stage1_col87[19] <= 1'b0;
                    stage1_col87[20] <= 1'b0;
                    stage1_col87[21] <= 1'b0;
                    stage1_col87[22] <= 1'b0;
                    stage1_col88[0] <= 1'b0;
                    stage1_col88[1] <= 1'b0;
                    stage1_col88[2] <= 1'b0;
                    stage1_col88[3] <= 1'b0;
                    stage1_col88[4] <= 1'b0;
                    stage1_col88[5] <= 1'b0;
                    stage1_col88[6] <= 1'b0;
                    stage1_col88[7] <= 1'b0;
                    stage1_col88[8] <= 1'b0;
                    stage1_col88[9] <= 1'b0;
                    stage1_col88[10] <= 1'b0;
                    stage1_col88[11] <= 1'b0;
                    stage1_col88[12] <= 1'b0;
                    stage1_col88[13] <= 1'b0;
                    stage1_col88[14] <= 1'b0;
                    stage1_col88[15] <= 1'b0;
                    stage1_col88[16] <= 1'b0;
                    stage1_col88[17] <= 1'b0;
                    stage1_col88[18] <= 1'b0;
                    stage1_col88[19] <= 1'b0;
                    stage1_col88[20] <= 1'b0;
                    stage1_col89[0] <= 1'b0;
                    stage1_col89[1] <= 1'b0;
                    stage1_col89[2] <= 1'b0;
                    stage1_col89[3] <= 1'b0;
                    stage1_col89[4] <= 1'b0;
                    stage1_col89[5] <= 1'b0;
                    stage1_col89[6] <= 1'b0;
                    stage1_col89[7] <= 1'b0;
                    stage1_col89[8] <= 1'b0;
                    stage1_col89[9] <= 1'b0;
                    stage1_col89[10] <= 1'b0;
                    stage1_col89[11] <= 1'b0;
                    stage1_col89[12] <= 1'b0;
                    stage1_col89[13] <= 1'b0;
                    stage1_col89[14] <= 1'b0;
                    stage1_col89[15] <= 1'b0;
                    stage1_col89[16] <= 1'b0;
                    stage1_col89[17] <= 1'b0;
                    stage1_col89[18] <= 1'b0;
                    stage1_col89[19] <= 1'b0;
                    stage1_col89[20] <= 1'b0;
                    stage1_col89[21] <= 1'b0;
                    stage1_col89[22] <= 1'b0;
                    stage1_col90[0] <= 1'b0;
                    stage1_col90[1] <= 1'b0;
                    stage1_col90[2] <= 1'b0;
                    stage1_col90[3] <= 1'b0;
                    stage1_col90[4] <= 1'b0;
                    stage1_col90[5] <= 1'b0;
                    stage1_col90[6] <= 1'b0;
                    stage1_col90[7] <= 1'b0;
                    stage1_col90[8] <= 1'b0;
                    stage1_col90[9] <= 1'b0;
                    stage1_col90[10] <= 1'b0;
                    stage1_col90[11] <= 1'b0;
                    stage1_col90[12] <= 1'b0;
                    stage1_col90[13] <= 1'b0;
                    stage1_col90[14] <= 1'b0;
                    stage1_col90[15] <= 1'b0;
                    stage1_col90[16] <= 1'b0;
                    stage1_col90[17] <= 1'b0;
                    stage1_col90[18] <= 1'b0;
                    stage1_col90[19] <= 1'b0;
                    stage1_col90[20] <= 1'b0;
                    stage1_col91[0] <= 1'b0;
                    stage1_col91[1] <= 1'b0;
                    stage1_col91[2] <= 1'b0;
                    stage1_col91[3] <= 1'b0;
                    stage1_col91[4] <= 1'b0;
                    stage1_col91[5] <= 1'b0;
                    stage1_col91[6] <= 1'b0;
                    stage1_col91[7] <= 1'b0;
                    stage1_col91[8] <= 1'b0;
                    stage1_col91[9] <= 1'b0;
                    stage1_col91[10] <= 1'b0;
                    stage1_col91[11] <= 1'b0;
                    stage1_col91[12] <= 1'b0;
                    stage1_col91[13] <= 1'b0;
                    stage1_col91[14] <= 1'b0;
                    stage1_col91[15] <= 1'b0;
                    stage1_col91[16] <= 1'b0;
                    stage1_col91[17] <= 1'b0;
                    stage1_col91[18] <= 1'b0;
                    stage1_col91[19] <= 1'b0;
                    stage1_col91[20] <= 1'b0;
                    stage1_col91[21] <= 1'b0;
                    stage1_col91[22] <= 1'b0;
                    stage1_col92[0] <= 1'b0;
                    stage1_col92[1] <= 1'b0;
                    stage1_col92[2] <= 1'b0;
                    stage1_col92[3] <= 1'b0;
                    stage1_col92[4] <= 1'b0;
                    stage1_col92[5] <= 1'b0;
                    stage1_col92[6] <= 1'b0;
                    stage1_col92[7] <= 1'b0;
                    stage1_col92[8] <= 1'b0;
                    stage1_col92[9] <= 1'b0;
                    stage1_col92[10] <= 1'b0;
                    stage1_col92[11] <= 1'b0;
                    stage1_col92[12] <= 1'b0;
                    stage1_col92[13] <= 1'b0;
                    stage1_col92[14] <= 1'b0;
                    stage1_col92[15] <= 1'b0;
                    stage1_col92[16] <= 1'b0;
                    stage1_col92[17] <= 1'b0;
                    stage1_col92[18] <= 1'b0;
                    stage1_col92[19] <= 1'b0;
                    stage1_col92[20] <= 1'b0;
                    stage1_col93[0] <= 1'b0;
                    stage1_col93[1] <= 1'b0;
                    stage1_col93[2] <= 1'b0;
                    stage1_col93[3] <= 1'b0;
                    stage1_col93[4] <= 1'b0;
                    stage1_col93[5] <= 1'b0;
                    stage1_col93[6] <= 1'b0;
                    stage1_col93[7] <= 1'b0;
                    stage1_col93[8] <= 1'b0;
                    stage1_col93[9] <= 1'b0;
                    stage1_col93[10] <= 1'b0;
                    stage1_col93[11] <= 1'b0;
                    stage1_col93[12] <= 1'b0;
                    stage1_col93[13] <= 1'b0;
                    stage1_col93[14] <= 1'b0;
                    stage1_col93[15] <= 1'b0;
                    stage1_col93[16] <= 1'b0;
                    stage1_col93[17] <= 1'b0;
                    stage1_col93[18] <= 1'b0;
                    stage1_col93[19] <= 1'b0;
                    stage1_col93[20] <= 1'b0;
                    stage1_col93[21] <= 1'b0;
                    stage1_col93[22] <= 1'b0;
                    stage1_col94[0] <= 1'b0;
                    stage1_col94[1] <= 1'b0;
                    stage1_col94[2] <= 1'b0;
                    stage1_col94[3] <= 1'b0;
                    stage1_col94[4] <= 1'b0;
                    stage1_col94[5] <= 1'b0;
                    stage1_col94[6] <= 1'b0;
                    stage1_col94[7] <= 1'b0;
                    stage1_col94[8] <= 1'b0;
                    stage1_col94[9] <= 1'b0;
                    stage1_col94[10] <= 1'b0;
                    stage1_col94[11] <= 1'b0;
                    stage1_col94[12] <= 1'b0;
                    stage1_col94[13] <= 1'b0;
                    stage1_col94[14] <= 1'b0;
                    stage1_col94[15] <= 1'b0;
                    stage1_col94[16] <= 1'b0;
                    stage1_col94[17] <= 1'b0;
                    stage1_col94[18] <= 1'b0;
                    stage1_col94[19] <= 1'b0;
                    stage1_col94[20] <= 1'b0;
                    stage1_col95[0] <= 1'b0;
                    stage1_col95[1] <= 1'b0;
                    stage1_col95[2] <= 1'b0;
                    stage1_col95[3] <= 1'b0;
                    stage1_col95[4] <= 1'b0;
                    stage1_col95[5] <= 1'b0;
                    stage1_col95[6] <= 1'b0;
                    stage1_col95[7] <= 1'b0;
                    stage1_col95[8] <= 1'b0;
                    stage1_col95[9] <= 1'b0;
                    stage1_col95[10] <= 1'b0;
                    stage1_col95[11] <= 1'b0;
                    stage1_col95[12] <= 1'b0;
                    stage1_col95[13] <= 1'b0;
                    stage1_col95[14] <= 1'b0;
                    stage1_col95[15] <= 1'b0;
                    stage1_col95[16] <= 1'b0;
                    stage1_col95[17] <= 1'b0;
                    stage1_col95[18] <= 1'b0;
                    stage1_col95[19] <= 1'b0;
                    stage1_col95[20] <= 1'b0;
                    stage1_col95[21] <= 1'b0;
                    stage1_col95[22] <= 1'b0;
                    stage1_col96[0] <= 1'b0;
                    stage1_col96[1] <= 1'b0;
                    stage1_col96[2] <= 1'b0;
                    stage1_col96[3] <= 1'b0;
                    stage1_col96[4] <= 1'b0;
                    stage1_col96[5] <= 1'b0;
                    stage1_col96[6] <= 1'b0;
                    stage1_col96[7] <= 1'b0;
                    stage1_col96[8] <= 1'b0;
                    stage1_col96[9] <= 1'b0;
                    stage1_col96[10] <= 1'b0;
                    stage1_col96[11] <= 1'b0;
                    stage1_col96[12] <= 1'b0;
                    stage1_col96[13] <= 1'b0;
                    stage1_col96[14] <= 1'b0;
                    stage1_col96[15] <= 1'b0;
                    stage1_col96[16] <= 1'b0;
                    stage1_col96[17] <= 1'b0;
                    stage1_col96[18] <= 1'b0;
                    stage1_col96[19] <= 1'b0;
                    stage1_col96[20] <= 1'b0;
                    stage1_col97[0] <= 1'b0;
                    stage1_col97[1] <= 1'b0;
                    stage1_col97[2] <= 1'b0;
                    stage1_col97[3] <= 1'b0;
                    stage1_col97[4] <= 1'b0;
                    stage1_col97[5] <= 1'b0;
                    stage1_col97[6] <= 1'b0;
                    stage1_col97[7] <= 1'b0;
                    stage1_col97[8] <= 1'b0;
                    stage1_col97[9] <= 1'b0;
                    stage1_col97[10] <= 1'b0;
                    stage1_col97[11] <= 1'b0;
                    stage1_col97[12] <= 1'b0;
                    stage1_col97[13] <= 1'b0;
                    stage1_col97[14] <= 1'b0;
                    stage1_col97[15] <= 1'b0;
                    stage1_col97[16] <= 1'b0;
                    stage1_col97[17] <= 1'b0;
                    stage1_col97[18] <= 1'b0;
                    stage1_col97[19] <= 1'b0;
                    stage1_col97[20] <= 1'b0;
                    stage1_col97[21] <= 1'b0;
                    stage1_col97[22] <= 1'b0;
                    stage1_col98[0] <= 1'b0;
                    stage1_col98[1] <= 1'b0;
                    stage1_col98[2] <= 1'b0;
                    stage1_col98[3] <= 1'b0;
                    stage1_col98[4] <= 1'b0;
                    stage1_col98[5] <= 1'b0;
                    stage1_col98[6] <= 1'b0;
                    stage1_col98[7] <= 1'b0;
                    stage1_col98[8] <= 1'b0;
                    stage1_col98[9] <= 1'b0;
                    stage1_col98[10] <= 1'b0;
                    stage1_col98[11] <= 1'b0;
                    stage1_col98[12] <= 1'b0;
                    stage1_col98[13] <= 1'b0;
                    stage1_col98[14] <= 1'b0;
                    stage1_col98[15] <= 1'b0;
                    stage1_col98[16] <= 1'b0;
                    stage1_col98[17] <= 1'b0;
                    stage1_col98[18] <= 1'b0;
                    stage1_col98[19] <= 1'b0;
                    stage1_col98[20] <= 1'b0;
                    stage1_col99[0] <= 1'b0;
                    stage1_col99[1] <= 1'b0;
                    stage1_col99[2] <= 1'b0;
                    stage1_col99[3] <= 1'b0;
                    stage1_col99[4] <= 1'b0;
                    stage1_col99[5] <= 1'b0;
                    stage1_col99[6] <= 1'b0;
                    stage1_col99[7] <= 1'b0;
                    stage1_col99[8] <= 1'b0;
                    stage1_col99[9] <= 1'b0;
                    stage1_col99[10] <= 1'b0;
                    stage1_col99[11] <= 1'b0;
                    stage1_col99[12] <= 1'b0;
                    stage1_col99[13] <= 1'b0;
                    stage1_col99[14] <= 1'b0;
                    stage1_col99[15] <= 1'b0;
                    stage1_col99[16] <= 1'b0;
                    stage1_col99[17] <= 1'b0;
                    stage1_col99[18] <= 1'b0;
                    stage1_col99[19] <= 1'b0;
                    stage1_col99[20] <= 1'b0;
                    stage1_col99[21] <= 1'b0;
                    stage1_col99[22] <= 1'b0;
                    stage1_col100[0] <= 1'b0;
                    stage1_col100[1] <= 1'b0;
                    stage1_col100[2] <= 1'b0;
                    stage1_col100[3] <= 1'b0;
                    stage1_col100[4] <= 1'b0;
                    stage1_col100[5] <= 1'b0;
                    stage1_col100[6] <= 1'b0;
                    stage1_col100[7] <= 1'b0;
                    stage1_col100[8] <= 1'b0;
                    stage1_col100[9] <= 1'b0;
                    stage1_col100[10] <= 1'b0;
                    stage1_col100[11] <= 1'b0;
                    stage1_col100[12] <= 1'b0;
                    stage1_col100[13] <= 1'b0;
                    stage1_col100[14] <= 1'b0;
                    stage1_col100[15] <= 1'b0;
                    stage1_col100[16] <= 1'b0;
                    stage1_col100[17] <= 1'b0;
                    stage1_col100[18] <= 1'b0;
                    stage1_col100[19] <= 1'b0;
                    stage1_col100[20] <= 1'b0;
                    stage1_col101[0] <= 1'b0;
                    stage1_col101[1] <= 1'b0;
                    stage1_col101[2] <= 1'b0;
                    stage1_col101[3] <= 1'b0;
                    stage1_col101[4] <= 1'b0;
                    stage1_col101[5] <= 1'b0;
                    stage1_col101[6] <= 1'b0;
                    stage1_col101[7] <= 1'b0;
                    stage1_col101[8] <= 1'b0;
                    stage1_col101[9] <= 1'b0;
                    stage1_col101[10] <= 1'b0;
                    stage1_col101[11] <= 1'b0;
                    stage1_col101[12] <= 1'b0;
                    stage1_col101[13] <= 1'b0;
                    stage1_col101[14] <= 1'b0;
                    stage1_col101[15] <= 1'b0;
                    stage1_col101[16] <= 1'b0;
                    stage1_col101[17] <= 1'b0;
                    stage1_col101[18] <= 1'b0;
                    stage1_col101[19] <= 1'b0;
                    stage1_col101[20] <= 1'b0;
                    stage1_col101[21] <= 1'b0;
                    stage1_col101[22] <= 1'b0;
                    stage1_col102[0] <= 1'b0;
                    stage1_col102[1] <= 1'b0;
                    stage1_col102[2] <= 1'b0;
                    stage1_col102[3] <= 1'b0;
                    stage1_col102[4] <= 1'b0;
                    stage1_col102[5] <= 1'b0;
                    stage1_col102[6] <= 1'b0;
                    stage1_col102[7] <= 1'b0;
                    stage1_col102[8] <= 1'b0;
                    stage1_col102[9] <= 1'b0;
                    stage1_col102[10] <= 1'b0;
                    stage1_col102[11] <= 1'b0;
                    stage1_col102[12] <= 1'b0;
                    stage1_col102[13] <= 1'b0;
                    stage1_col102[14] <= 1'b0;
                    stage1_col102[15] <= 1'b0;
                    stage1_col102[16] <= 1'b0;
                    stage1_col102[17] <= 1'b0;
                    stage1_col102[18] <= 1'b0;
                    stage1_col102[19] <= 1'b0;
                    stage1_col102[20] <= 1'b0;
                    stage1_col103[0] <= 1'b0;
                    stage1_col103[1] <= 1'b0;
                    stage1_col103[2] <= 1'b0;
                    stage1_col103[3] <= 1'b0;
                    stage1_col103[4] <= 1'b0;
                    stage1_col103[5] <= 1'b0;
                    stage1_col103[6] <= 1'b0;
                    stage1_col103[7] <= 1'b0;
                    stage1_col103[8] <= 1'b0;
                    stage1_col103[9] <= 1'b0;
                    stage1_col103[10] <= 1'b0;
                    stage1_col103[11] <= 1'b0;
                    stage1_col103[12] <= 1'b0;
                    stage1_col103[13] <= 1'b0;
                    stage1_col103[14] <= 1'b0;
                    stage1_col103[15] <= 1'b0;
                    stage1_col103[16] <= 1'b0;
                    stage1_col103[17] <= 1'b0;
                    stage1_col103[18] <= 1'b0;
                    stage1_col103[19] <= 1'b0;
                    stage1_col103[20] <= 1'b0;
                    stage1_col103[21] <= 1'b0;
                    stage1_col103[22] <= 1'b0;
                    stage1_col104[0] <= 1'b0;
                    stage1_col104[1] <= 1'b0;
                    stage1_col104[2] <= 1'b0;
                    stage1_col104[3] <= 1'b0;
                    stage1_col104[4] <= 1'b0;
                    stage1_col104[5] <= 1'b0;
                    stage1_col104[6] <= 1'b0;
                    stage1_col104[7] <= 1'b0;
                    stage1_col104[8] <= 1'b0;
                    stage1_col104[9] <= 1'b0;
                    stage1_col104[10] <= 1'b0;
                    stage1_col104[11] <= 1'b0;
                    stage1_col104[12] <= 1'b0;
                    stage1_col104[13] <= 1'b0;
                    stage1_col104[14] <= 1'b0;
                    stage1_col104[15] <= 1'b0;
                    stage1_col104[16] <= 1'b0;
                    stage1_col104[17] <= 1'b0;
                    stage1_col104[18] <= 1'b0;
                    stage1_col104[19] <= 1'b0;
                    stage1_col104[20] <= 1'b0;
                    stage1_col105[0] <= 1'b0;
                    stage1_col105[1] <= 1'b0;
                    stage1_col105[2] <= 1'b0;
                    stage1_col105[3] <= 1'b0;
                    stage1_col105[4] <= 1'b0;
                    stage1_col105[5] <= 1'b0;
                    stage1_col105[6] <= 1'b0;
                    stage1_col105[7] <= 1'b0;
                    stage1_col105[8] <= 1'b0;
                    stage1_col105[9] <= 1'b0;
                    stage1_col105[10] <= 1'b0;
                    stage1_col105[11] <= 1'b0;
                    stage1_col105[12] <= 1'b0;
                    stage1_col105[13] <= 1'b0;
                    stage1_col105[14] <= 1'b0;
                    stage1_col105[15] <= 1'b0;
                    stage1_col105[16] <= 1'b0;
                    stage1_col105[17] <= 1'b0;
                    stage1_col105[18] <= 1'b0;
                    stage1_col105[19] <= 1'b0;
                    stage1_col105[20] <= 1'b0;
                    stage1_col105[21] <= 1'b0;
                    stage1_col105[22] <= 1'b0;
                    stage1_col106[0] <= 1'b0;
                    stage1_col106[1] <= 1'b0;
                    stage1_col106[2] <= 1'b0;
                    stage1_col106[3] <= 1'b0;
                    stage1_col106[4] <= 1'b0;
                    stage1_col106[5] <= 1'b0;
                    stage1_col106[6] <= 1'b0;
                    stage1_col106[7] <= 1'b0;
                    stage1_col106[8] <= 1'b0;
                    stage1_col106[9] <= 1'b0;
                    stage1_col106[10] <= 1'b0;
                    stage1_col106[11] <= 1'b0;
                    stage1_col106[12] <= 1'b0;
                    stage1_col106[13] <= 1'b0;
                    stage1_col106[14] <= 1'b0;
                    stage1_col106[15] <= 1'b0;
                    stage1_col106[16] <= 1'b0;
                    stage1_col106[17] <= 1'b0;
                    stage1_col106[18] <= 1'b0;
                    stage1_col106[19] <= 1'b0;
                    stage1_col106[20] <= 1'b0;
                    stage1_col107[0] <= 1'b0;
                    stage1_col107[1] <= 1'b0;
                    stage1_col107[2] <= 1'b0;
                    stage1_col107[3] <= 1'b0;
                    stage1_col107[4] <= 1'b0;
                    stage1_col107[5] <= 1'b0;
                    stage1_col107[6] <= 1'b0;
                    stage1_col107[7] <= 1'b0;
                    stage1_col107[8] <= 1'b0;
                    stage1_col107[9] <= 1'b0;
                    stage1_col107[10] <= 1'b0;
                    stage1_col107[11] <= 1'b0;
                    stage1_col107[12] <= 1'b0;
                    stage1_col107[13] <= 1'b0;
                    stage1_col107[14] <= 1'b0;
                    stage1_col107[15] <= 1'b0;
                    stage1_col107[16] <= 1'b0;
                    stage1_col107[17] <= 1'b0;
                    stage1_col107[18] <= 1'b0;
                    stage1_col107[19] <= 1'b0;
                    stage1_col107[20] <= 1'b0;
                    stage1_col107[21] <= 1'b0;
                    stage1_col107[22] <= 1'b0;
                    stage1_col108[0] <= 1'b0;
                    stage1_col108[1] <= 1'b0;
                    stage1_col108[2] <= 1'b0;
                    stage1_col108[3] <= 1'b0;
                    stage1_col108[4] <= 1'b0;
                    stage1_col108[5] <= 1'b0;
                    stage1_col108[6] <= 1'b0;
                    stage1_col108[7] <= 1'b0;
                    stage1_col108[8] <= 1'b0;
                    stage1_col108[9] <= 1'b0;
                    stage1_col108[10] <= 1'b0;
                    stage1_col108[11] <= 1'b0;
                    stage1_col108[12] <= 1'b0;
                    stage1_col108[13] <= 1'b0;
                    stage1_col108[14] <= 1'b0;
                    stage1_col108[15] <= 1'b0;
                    stage1_col108[16] <= 1'b0;
                    stage1_col108[17] <= 1'b0;
                    stage1_col108[18] <= 1'b0;
                    stage1_col108[19] <= 1'b0;
                    stage1_col108[20] <= 1'b0;
                    stage1_col109[0] <= 1'b0;
                    stage1_col109[1] <= 1'b0;
                    stage1_col109[2] <= 1'b0;
                    stage1_col109[3] <= 1'b0;
                    stage1_col109[4] <= 1'b0;
                    stage1_col109[5] <= 1'b0;
                    stage1_col109[6] <= 1'b0;
                    stage1_col109[7] <= 1'b0;
                    stage1_col109[8] <= 1'b0;
                    stage1_col109[9] <= 1'b0;
                    stage1_col109[10] <= 1'b0;
                    stage1_col109[11] <= 1'b0;
                    stage1_col109[12] <= 1'b0;
                    stage1_col109[13] <= 1'b0;
                    stage1_col109[14] <= 1'b0;
                    stage1_col109[15] <= 1'b0;
                    stage1_col109[16] <= 1'b0;
                    stage1_col109[17] <= 1'b0;
                    stage1_col109[18] <= 1'b0;
                    stage1_col109[19] <= 1'b0;
                    stage1_col109[20] <= 1'b0;
                    stage1_col109[21] <= 1'b0;
                    stage1_col109[22] <= 1'b0;
                    stage1_col110[0] <= 1'b0;
                    stage1_col110[1] <= 1'b0;
                    stage1_col110[2] <= 1'b0;
                    stage1_col110[3] <= 1'b0;
                    stage1_col110[4] <= 1'b0;
                    stage1_col110[5] <= 1'b0;
                    stage1_col110[6] <= 1'b0;
                    stage1_col110[7] <= 1'b0;
                    stage1_col110[8] <= 1'b0;
                    stage1_col110[9] <= 1'b0;
                    stage1_col110[10] <= 1'b0;
                    stage1_col110[11] <= 1'b0;
                    stage1_col110[12] <= 1'b0;
                    stage1_col110[13] <= 1'b0;
                    stage1_col110[14] <= 1'b0;
                    stage1_col110[15] <= 1'b0;
                    stage1_col110[16] <= 1'b0;
                    stage1_col110[17] <= 1'b0;
                    stage1_col110[18] <= 1'b0;
                    stage1_col110[19] <= 1'b0;
                    stage1_col110[20] <= 1'b0;
                    stage1_col111[0] <= 1'b0;
                    stage1_col111[1] <= 1'b0;
                    stage1_col111[2] <= 1'b0;
                    stage1_col111[3] <= 1'b0;
                    stage1_col111[4] <= 1'b0;
                    stage1_col111[5] <= 1'b0;
                    stage1_col111[6] <= 1'b0;
                    stage1_col111[7] <= 1'b0;
                    stage1_col111[8] <= 1'b0;
                    stage1_col111[9] <= 1'b0;
                    stage1_col111[10] <= 1'b0;
                    stage1_col111[11] <= 1'b0;
                    stage1_col111[12] <= 1'b0;
                    stage1_col111[13] <= 1'b0;
                    stage1_col111[14] <= 1'b0;
                    stage1_col111[15] <= 1'b0;
                    stage1_col111[16] <= 1'b0;
                    stage1_col111[17] <= 1'b0;
                    stage1_col111[18] <= 1'b0;
                    stage1_col111[19] <= 1'b0;
                    stage1_col111[20] <= 1'b0;
                    stage1_col111[21] <= 1'b0;
                    stage1_col111[22] <= 1'b0;
                    stage1_col112[0] <= 1'b0;
                    stage1_col112[1] <= 1'b0;
                    stage1_col112[2] <= 1'b0;
                    stage1_col112[3] <= 1'b0;
                    stage1_col112[4] <= 1'b0;
                    stage1_col112[5] <= 1'b0;
                    stage1_col112[6] <= 1'b0;
                    stage1_col112[7] <= 1'b0;
                    stage1_col112[8] <= 1'b0;
                    stage1_col112[9] <= 1'b0;
                    stage1_col112[10] <= 1'b0;
                    stage1_col112[11] <= 1'b0;
                    stage1_col112[12] <= 1'b0;
                    stage1_col112[13] <= 1'b0;
                    stage1_col112[14] <= 1'b0;
                    stage1_col112[15] <= 1'b0;
                    stage1_col112[16] <= 1'b0;
                    stage1_col112[17] <= 1'b0;
                    stage1_col112[18] <= 1'b0;
                    stage1_col112[19] <= 1'b0;
                    stage1_col112[20] <= 1'b0;
                    stage1_col113[0] <= 1'b0;
                    stage1_col113[1] <= 1'b0;
                    stage1_col113[2] <= 1'b0;
                    stage1_col113[3] <= 1'b0;
                    stage1_col113[4] <= 1'b0;
                    stage1_col113[5] <= 1'b0;
                    stage1_col113[6] <= 1'b0;
                    stage1_col113[7] <= 1'b0;
                    stage1_col113[8] <= 1'b0;
                    stage1_col113[9] <= 1'b0;
                    stage1_col113[10] <= 1'b0;
                    stage1_col113[11] <= 1'b0;
                    stage1_col113[12] <= 1'b0;
                    stage1_col113[13] <= 1'b0;
                    stage1_col113[14] <= 1'b0;
                    stage1_col113[15] <= 1'b0;
                    stage1_col113[16] <= 1'b0;
                    stage1_col113[17] <= 1'b0;
                    stage1_col113[18] <= 1'b0;
                    stage1_col113[19] <= 1'b0;
                    stage1_col113[20] <= 1'b0;
                    stage1_col113[21] <= 1'b0;
                    stage1_col113[22] <= 1'b0;
                    stage1_col114[0] <= 1'b0;
                    stage1_col114[1] <= 1'b0;
                    stage1_col114[2] <= 1'b0;
                    stage1_col114[3] <= 1'b0;
                    stage1_col114[4] <= 1'b0;
                    stage1_col114[5] <= 1'b0;
                    stage1_col114[6] <= 1'b0;
                    stage1_col114[7] <= 1'b0;
                    stage1_col114[8] <= 1'b0;
                    stage1_col114[9] <= 1'b0;
                    stage1_col114[10] <= 1'b0;
                    stage1_col114[11] <= 1'b0;
                    stage1_col114[12] <= 1'b0;
                    stage1_col114[13] <= 1'b0;
                    stage1_col114[14] <= 1'b0;
                    stage1_col114[15] <= 1'b0;
                    stage1_col114[16] <= 1'b0;
                    stage1_col114[17] <= 1'b0;
                    stage1_col114[18] <= 1'b0;
                    stage1_col114[19] <= 1'b0;
                    stage1_col114[20] <= 1'b0;
                    stage1_col115[0] <= 1'b0;
                    stage1_col115[1] <= 1'b0;
                    stage1_col115[2] <= 1'b0;
                    stage1_col115[3] <= 1'b0;
                    stage1_col115[4] <= 1'b0;
                    stage1_col115[5] <= 1'b0;
                    stage1_col115[6] <= 1'b0;
                    stage1_col115[7] <= 1'b0;
                    stage1_col115[8] <= 1'b0;
                    stage1_col115[9] <= 1'b0;
                    stage1_col115[10] <= 1'b0;
                    stage1_col115[11] <= 1'b0;
                    stage1_col115[12] <= 1'b0;
                    stage1_col115[13] <= 1'b0;
                    stage1_col115[14] <= 1'b0;
                    stage1_col115[15] <= 1'b0;
                    stage1_col115[16] <= 1'b0;
                    stage1_col115[17] <= 1'b0;
                    stage1_col115[18] <= 1'b0;
                    stage1_col115[19] <= 1'b0;
                    stage1_col115[20] <= 1'b0;
                    stage1_col115[21] <= 1'b0;
                    stage1_col115[22] <= 1'b0;
                    stage1_col116[0] <= 1'b0;
                    stage1_col116[1] <= 1'b0;
                    stage1_col116[2] <= 1'b0;
                    stage1_col116[3] <= 1'b0;
                    stage1_col116[4] <= 1'b0;
                    stage1_col116[5] <= 1'b0;
                    stage1_col116[6] <= 1'b0;
                    stage1_col116[7] <= 1'b0;
                    stage1_col116[8] <= 1'b0;
                    stage1_col116[9] <= 1'b0;
                    stage1_col116[10] <= 1'b0;
                    stage1_col116[11] <= 1'b0;
                    stage1_col116[12] <= 1'b0;
                    stage1_col116[13] <= 1'b0;
                    stage1_col116[14] <= 1'b0;
                    stage1_col116[15] <= 1'b0;
                    stage1_col116[16] <= 1'b0;
                    stage1_col116[17] <= 1'b0;
                    stage1_col116[18] <= 1'b0;
                    stage1_col116[19] <= 1'b0;
                    stage1_col116[20] <= 1'b0;
                    stage1_col117[0] <= 1'b0;
                    stage1_col117[1] <= 1'b0;
                    stage1_col117[2] <= 1'b0;
                    stage1_col117[3] <= 1'b0;
                    stage1_col117[4] <= 1'b0;
                    stage1_col117[5] <= 1'b0;
                    stage1_col117[6] <= 1'b0;
                    stage1_col117[7] <= 1'b0;
                    stage1_col117[8] <= 1'b0;
                    stage1_col117[9] <= 1'b0;
                    stage1_col117[10] <= 1'b0;
                    stage1_col117[11] <= 1'b0;
                    stage1_col117[12] <= 1'b0;
                    stage1_col117[13] <= 1'b0;
                    stage1_col117[14] <= 1'b0;
                    stage1_col117[15] <= 1'b0;
                    stage1_col117[16] <= 1'b0;
                    stage1_col117[17] <= 1'b0;
                    stage1_col117[18] <= 1'b0;
                    stage1_col117[19] <= 1'b0;
                    stage1_col117[20] <= 1'b0;
                    stage1_col117[21] <= 1'b0;
                    stage1_col117[22] <= 1'b0;
                    stage1_col118[0] <= 1'b0;
                    stage1_col118[1] <= 1'b0;
                    stage1_col118[2] <= 1'b0;
                    stage1_col118[3] <= 1'b0;
                    stage1_col118[4] <= 1'b0;
                    stage1_col118[5] <= 1'b0;
                    stage1_col118[6] <= 1'b0;
                    stage1_col118[7] <= 1'b0;
                    stage1_col118[8] <= 1'b0;
                    stage1_col118[9] <= 1'b0;
                    stage1_col118[10] <= 1'b0;
                    stage1_col118[11] <= 1'b0;
                    stage1_col118[12] <= 1'b0;
                    stage1_col118[13] <= 1'b0;
                    stage1_col118[14] <= 1'b0;
                    stage1_col118[15] <= 1'b0;
                    stage1_col118[16] <= 1'b0;
                    stage1_col118[17] <= 1'b0;
                    stage1_col118[18] <= 1'b0;
                    stage1_col118[19] <= 1'b0;
                    stage1_col118[20] <= 1'b0;
                    stage1_col119[0] <= 1'b0;
                    stage1_col119[1] <= 1'b0;
                    stage1_col119[2] <= 1'b0;
                    stage1_col119[3] <= 1'b0;
                    stage1_col119[4] <= 1'b0;
                    stage1_col119[5] <= 1'b0;
                    stage1_col119[6] <= 1'b0;
                    stage1_col119[7] <= 1'b0;
                    stage1_col119[8] <= 1'b0;
                    stage1_col119[9] <= 1'b0;
                    stage1_col119[10] <= 1'b0;
                    stage1_col119[11] <= 1'b0;
                    stage1_col119[12] <= 1'b0;
                    stage1_col119[13] <= 1'b0;
                    stage1_col119[14] <= 1'b0;
                    stage1_col119[15] <= 1'b0;
                    stage1_col119[16] <= 1'b0;
                    stage1_col119[17] <= 1'b0;
                    stage1_col119[18] <= 1'b0;
                    stage1_col119[19] <= 1'b0;
                    stage1_col119[20] <= 1'b0;
                    stage1_col119[21] <= 1'b0;
                    stage1_col119[22] <= 1'b0;
                    stage1_col120[0] <= 1'b0;
                    stage1_col120[1] <= 1'b0;
                    stage1_col120[2] <= 1'b0;
                    stage1_col120[3] <= 1'b0;
                    stage1_col120[4] <= 1'b0;
                    stage1_col120[5] <= 1'b0;
                    stage1_col120[6] <= 1'b0;
                    stage1_col120[7] <= 1'b0;
                    stage1_col120[8] <= 1'b0;
                    stage1_col120[9] <= 1'b0;
                    stage1_col120[10] <= 1'b0;
                    stage1_col120[11] <= 1'b0;
                    stage1_col120[12] <= 1'b0;
                    stage1_col120[13] <= 1'b0;
                    stage1_col120[14] <= 1'b0;
                    stage1_col120[15] <= 1'b0;
                    stage1_col120[16] <= 1'b0;
                    stage1_col120[17] <= 1'b0;
                    stage1_col120[18] <= 1'b0;
                    stage1_col120[19] <= 1'b0;
                    stage1_col120[20] <= 1'b0;
                    stage1_col121[0] <= 1'b0;
                    stage1_col121[1] <= 1'b0;
                    stage1_col121[2] <= 1'b0;
                    stage1_col121[3] <= 1'b0;
                    stage1_col121[4] <= 1'b0;
                    stage1_col121[5] <= 1'b0;
                    stage1_col121[6] <= 1'b0;
                    stage1_col121[7] <= 1'b0;
                    stage1_col121[8] <= 1'b0;
                    stage1_col121[9] <= 1'b0;
                    stage1_col121[10] <= 1'b0;
                    stage1_col121[11] <= 1'b0;
                    stage1_col121[12] <= 1'b0;
                    stage1_col121[13] <= 1'b0;
                    stage1_col121[14] <= 1'b0;
                    stage1_col121[15] <= 1'b0;
                    stage1_col121[16] <= 1'b0;
                    stage1_col121[17] <= 1'b0;
                    stage1_col121[18] <= 1'b0;
                    stage1_col121[19] <= 1'b0;
                    stage1_col121[20] <= 1'b0;
                    stage1_col121[21] <= 1'b0;
                    stage1_col121[22] <= 1'b0;
                    stage1_col122[0] <= 1'b0;
                    stage1_col122[1] <= 1'b0;
                    stage1_col122[2] <= 1'b0;
                    stage1_col122[3] <= 1'b0;
                    stage1_col122[4] <= 1'b0;
                    stage1_col122[5] <= 1'b0;
                    stage1_col122[6] <= 1'b0;
                    stage1_col122[7] <= 1'b0;
                    stage1_col122[8] <= 1'b0;
                    stage1_col122[9] <= 1'b0;
                    stage1_col122[10] <= 1'b0;
                    stage1_col122[11] <= 1'b0;
                    stage1_col122[12] <= 1'b0;
                    stage1_col122[13] <= 1'b0;
                    stage1_col122[14] <= 1'b0;
                    stage1_col122[15] <= 1'b0;
                    stage1_col122[16] <= 1'b0;
                    stage1_col122[17] <= 1'b0;
                    stage1_col122[18] <= 1'b0;
                    stage1_col122[19] <= 1'b0;
                    stage1_col122[20] <= 1'b0;
                    stage1_col123[0] <= 1'b0;
                    stage1_col123[1] <= 1'b0;
                    stage1_col123[2] <= 1'b0;
                    stage1_col123[3] <= 1'b0;
                    stage1_col123[4] <= 1'b0;
                    stage1_col123[5] <= 1'b0;
                    stage1_col123[6] <= 1'b0;
                    stage1_col123[7] <= 1'b0;
                    stage1_col123[8] <= 1'b0;
                    stage1_col123[9] <= 1'b0;
                    stage1_col123[10] <= 1'b0;
                    stage1_col123[11] <= 1'b0;
                    stage1_col123[12] <= 1'b0;
                    stage1_col123[13] <= 1'b0;
                    stage1_col123[14] <= 1'b0;
                    stage1_col123[15] <= 1'b0;
                    stage1_col123[16] <= 1'b0;
                    stage1_col123[17] <= 1'b0;
                    stage1_col123[18] <= 1'b0;
                    stage1_col123[19] <= 1'b0;
                    stage1_col123[20] <= 1'b0;
                    stage1_col123[21] <= 1'b0;
                    stage1_col123[22] <= 1'b0;
                    stage1_col124[0] <= 1'b0;
                    stage1_col124[1] <= 1'b0;
                    stage1_col124[2] <= 1'b0;
                    stage1_col124[3] <= 1'b0;
                    stage1_col124[4] <= 1'b0;
                    stage1_col124[5] <= 1'b0;
                    stage1_col124[6] <= 1'b0;
                    stage1_col124[7] <= 1'b0;
                    stage1_col124[8] <= 1'b0;
                    stage1_col124[9] <= 1'b0;
                    stage1_col124[10] <= 1'b0;
                    stage1_col124[11] <= 1'b0;
                    stage1_col124[12] <= 1'b0;
                    stage1_col124[13] <= 1'b0;
                    stage1_col124[14] <= 1'b0;
                    stage1_col124[15] <= 1'b0;
                    stage1_col124[16] <= 1'b0;
                    stage1_col124[17] <= 1'b0;
                    stage1_col124[18] <= 1'b0;
                    stage1_col124[19] <= 1'b0;
                    stage1_col124[20] <= 1'b0;
                    stage1_col125[0] <= 1'b0;
                    stage1_col125[1] <= 1'b0;
                    stage1_col125[2] <= 1'b0;
                    stage1_col125[3] <= 1'b0;
                    stage1_col125[4] <= 1'b0;
                    stage1_col125[5] <= 1'b0;
                    stage1_col125[6] <= 1'b0;
                    stage1_col125[7] <= 1'b0;
                    stage1_col125[8] <= 1'b0;
                    stage1_col125[9] <= 1'b0;
                    stage1_col125[10] <= 1'b0;
                    stage1_col125[11] <= 1'b0;
                    stage1_col125[12] <= 1'b0;
                    stage1_col125[13] <= 1'b0;
                    stage1_col125[14] <= 1'b0;
                    stage1_col125[15] <= 1'b0;
                    stage1_col125[16] <= 1'b0;
                    stage1_col125[17] <= 1'b0;
                    stage1_col125[18] <= 1'b0;
                    stage1_col125[19] <= 1'b0;
                    stage1_col125[20] <= 1'b0;
                    stage1_col125[21] <= 1'b0;
                    stage1_col125[22] <= 1'b0;
                    stage1_col126[0] <= 1'b0;
                    stage1_col126[1] <= 1'b0;
                    stage1_col126[2] <= 1'b0;
                    stage1_col126[3] <= 1'b0;
                    stage1_col126[4] <= 1'b0;
                    stage1_col126[5] <= 1'b0;
                    stage1_col126[6] <= 1'b0;
                    stage1_col126[7] <= 1'b0;
                    stage1_col126[8] <= 1'b0;
                    stage1_col126[9] <= 1'b0;
                    stage1_col126[10] <= 1'b0;
                    stage1_col126[11] <= 1'b0;
                    stage1_col126[12] <= 1'b0;
                    stage1_col126[13] <= 1'b0;
                    stage1_col126[14] <= 1'b0;
                    stage1_col126[15] <= 1'b0;
                    stage1_col126[16] <= 1'b0;
                    stage1_col126[17] <= 1'b0;
                    stage1_col126[18] <= 1'b0;
                    stage1_col126[19] <= 1'b0;
                    stage1_col126[20] <= 1'b0;
                    stage1_col127[0] <= 1'b0;
                    stage1_col127[1] <= 1'b0;
                    stage1_col127[2] <= 1'b0;
                    stage1_col127[3] <= 1'b0;
                    stage1_col127[4] <= 1'b0;
                    stage1_col127[5] <= 1'b0;
                    stage1_col127[6] <= 1'b0;
                    stage1_col127[7] <= 1'b0;
                    stage1_col127[8] <= 1'b0;
                    stage1_col127[9] <= 1'b0;
                    stage1_col127[10] <= 1'b0;
                    stage1_col127[11] <= 1'b0;
                    stage1_col127[12] <= 1'b0;
                    stage1_col127[13] <= 1'b0;
                    stage1_col127[14] <= 1'b0;
                    stage1_col127[15] <= 1'b0;
                    stage1_col127[16] <= 1'b0;
                    stage1_col127[17] <= 1'b0;
                    stage1_col127[18] <= 1'b0;
                    stage1_col127[19] <= 1'b0;
                    stage1_col127[20] <= 1'b0;
                    stage1_col127[21] <= 1'b0;
                    stage1_col127[22] <= 1'b0;
                    stage1_col127[23] <= 1'b0;
                    stage1_col127[24] <= 1'b0;
                    stage1_col127[25] <= 1'b0;
                    stage1_col127[26] <= 1'b0;
                    stage1_col127[27] <= 1'b0;
                    stage1_col127[28] <= 1'b0;
                    stage1_col127[29] <= 1'b0;
                    stage1_col127[30] <= 1'b0;
                    stage1_col127[31] <= 1'b0;
                    stage1_col127[32] <= 1'b0;
                    stage1_col127[33] <= 1'b0;
                    stage1_col127[34] <= 1'b0;
                    stage1_col127[35] <= 1'b0;
                    stage1_col127[36] <= 1'b0;
                    stage1_col127[37] <= 1'b0;
                    stage1_col127[38] <= 1'b0;
                    stage1_col127[39] <= 1'b0;
                    stage1_col127[40] <= 1'b0;
                    stage1_col127[41] <= 1'b0;
                    stage1_col127[42] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage1_col0[0] <= ha_s0_c0_n0_s;
                    stage1_col1[0] <= ha_s0_c0_n0_c;
                    stage1_col1[1] <= stage0_col1[0];
                    stage1_col2[0] <= fa_s0_c2_n0_s;
                    stage1_col3[0] <= fa_s0_c2_n0_c;
                    stage1_col3[1] <= stage0_col3[0];
                    stage1_col3[2] <= stage0_col3[1];
                    stage1_col4[0] <= fa_s0_c4_n1_s;
                    stage1_col4[1] <= stage0_col4[3];
                    stage1_col5[0] <= fa_s0_c4_n1_c;
                    stage1_col5[1] <= fa_s0_c5_n2_s;
                    stage1_col6[0] <= fa_s0_c5_n2_c;
                    stage1_col6[1] <= fa_s0_c6_n3_s;
                    stage1_col6[2] <= stage0_col6[3];
                    stage1_col6[3] <= stage0_col6[4];
                    stage1_col7[0] <= fa_s0_c6_n3_c;
                    stage1_col7[1] <= fa_s0_c7_n4_s;
                    stage1_col7[2] <= stage0_col7[3];
                    stage1_col8[0] <= fa_s0_c7_n4_c;
                    stage1_col8[1] <= fa_s0_c8_n5_s;
                    stage1_col8[2] <= fa_s0_c8_n6_s;
                    stage1_col9[0] <= fa_s0_c8_n5_c;
                    stage1_col9[1] <= fa_s0_c8_n6_c;
                    stage1_col9[2] <= fa_s0_c9_n7_s;
                    stage1_col9[3] <= stage0_col9[3];
                    stage1_col9[4] <= stage0_col9[4];
                    stage1_col10[0] <= fa_s0_c9_n7_c;
                    stage1_col10[1] <= fa_s0_c10_n8_s;
                    stage1_col10[2] <= fa_s0_c10_n9_s;
                    stage1_col10[3] <= stage0_col10[6];
                    stage1_col11[0] <= fa_s0_c10_n8_c;
                    stage1_col11[1] <= fa_s0_c10_n9_c;
                    stage1_col11[2] <= fa_s0_c11_n10_s;
                    stage1_col11[3] <= fa_s0_c11_n11_s;
                    stage1_col12[0] <= fa_s0_c11_n10_c;
                    stage1_col12[1] <= fa_s0_c11_n11_c;
                    stage1_col12[2] <= fa_s0_c12_n12_s;
                    stage1_col12[3] <= fa_s0_c12_n13_s;
                    stage1_col12[4] <= stage0_col12[6];
                    stage1_col12[5] <= stage0_col12[7];
                    stage1_col13[0] <= fa_s0_c12_n12_c;
                    stage1_col13[1] <= fa_s0_c12_n13_c;
                    stage1_col13[2] <= fa_s0_c13_n14_s;
                    stage1_col13[3] <= fa_s0_c13_n15_s;
                    stage1_col13[4] <= stage0_col13[6];
                    stage1_col14[0] <= fa_s0_c13_n14_c;
                    stage1_col14[1] <= fa_s0_c13_n15_c;
                    stage1_col14[2] <= fa_s0_c14_n16_s;
                    stage1_col14[3] <= fa_s0_c14_n17_s;
                    stage1_col14[4] <= fa_s0_c14_n18_s;
                    stage1_col15[0] <= fa_s0_c14_n16_c;
                    stage1_col15[1] <= fa_s0_c14_n17_c;
                    stage1_col15[2] <= fa_s0_c14_n18_c;
                    stage1_col15[3] <= fa_s0_c15_n19_s;
                    stage1_col15[4] <= fa_s0_c15_n20_s;
                    stage1_col15[5] <= stage0_col15[6];
                    stage1_col15[6] <= stage0_col15[7];
                    stage1_col16[0] <= fa_s0_c15_n19_c;
                    stage1_col16[1] <= fa_s0_c15_n20_c;
                    stage1_col16[2] <= fa_s0_c16_n21_s;
                    stage1_col16[3] <= fa_s0_c16_n22_s;
                    stage1_col16[4] <= fa_s0_c16_n23_s;
                    stage1_col16[5] <= stage0_col16[9];
                    stage1_col17[0] <= fa_s0_c16_n21_c;
                    stage1_col17[1] <= fa_s0_c16_n22_c;
                    stage1_col17[2] <= fa_s0_c16_n23_c;
                    stage1_col17[3] <= fa_s0_c17_n24_s;
                    stage1_col17[4] <= fa_s0_c17_n25_s;
                    stage1_col17[5] <= fa_s0_c17_n26_s;
                    stage1_col18[0] <= fa_s0_c17_n24_c;
                    stage1_col18[1] <= fa_s0_c17_n25_c;
                    stage1_col18[2] <= fa_s0_c17_n26_c;
                    stage1_col18[3] <= fa_s0_c18_n27_s;
                    stage1_col18[4] <= fa_s0_c18_n28_s;
                    stage1_col18[5] <= fa_s0_c18_n29_s;
                    stage1_col18[6] <= stage0_col18[9];
                    stage1_col18[7] <= stage0_col18[10];
                    stage1_col19[0] <= fa_s0_c18_n27_c;
                    stage1_col19[1] <= fa_s0_c18_n28_c;
                    stage1_col19[2] <= fa_s0_c18_n29_c;
                    stage1_col19[3] <= fa_s0_c19_n30_s;
                    stage1_col19[4] <= fa_s0_c19_n31_s;
                    stage1_col19[5] <= fa_s0_c19_n32_s;
                    stage1_col19[6] <= stage0_col19[9];
                    stage1_col20[0] <= fa_s0_c19_n30_c;
                    stage1_col20[1] <= fa_s0_c19_n31_c;
                    stage1_col20[2] <= fa_s0_c19_n32_c;
                    stage1_col20[3] <= fa_s0_c20_n33_s;
                    stage1_col20[4] <= fa_s0_c20_n34_s;
                    stage1_col20[5] <= fa_s0_c20_n35_s;
                    stage1_col20[6] <= fa_s0_c20_n36_s;
                    stage1_col21[0] <= fa_s0_c20_n33_c;
                    stage1_col21[1] <= fa_s0_c20_n34_c;
                    stage1_col21[2] <= fa_s0_c20_n35_c;
                    stage1_col21[3] <= fa_s0_c20_n36_c;
                    stage1_col21[4] <= fa_s0_c21_n37_s;
                    stage1_col21[5] <= fa_s0_c21_n38_s;
                    stage1_col21[6] <= fa_s0_c21_n39_s;
                    stage1_col21[7] <= stage0_col21[9];
                    stage1_col21[8] <= stage0_col21[10];
                    stage1_col22[0] <= fa_s0_c21_n37_c;
                    stage1_col22[1] <= fa_s0_c21_n38_c;
                    stage1_col22[2] <= fa_s0_c21_n39_c;
                    stage1_col22[3] <= fa_s0_c22_n40_s;
                    stage1_col22[4] <= fa_s0_c22_n41_s;
                    stage1_col22[5] <= fa_s0_c22_n42_s;
                    stage1_col22[6] <= fa_s0_c22_n43_s;
                    stage1_col22[7] <= stage0_col22[12];
                    stage1_col23[0] <= fa_s0_c22_n40_c;
                    stage1_col23[1] <= fa_s0_c22_n41_c;
                    stage1_col23[2] <= fa_s0_c22_n42_c;
                    stage1_col23[3] <= fa_s0_c22_n43_c;
                    stage1_col23[4] <= fa_s0_c23_n44_s;
                    stage1_col23[5] <= fa_s0_c23_n45_s;
                    stage1_col23[6] <= fa_s0_c23_n46_s;
                    stage1_col23[7] <= fa_s0_c23_n47_s;
                    stage1_col24[0] <= fa_s0_c23_n44_c;
                    stage1_col24[1] <= fa_s0_c23_n45_c;
                    stage1_col24[2] <= fa_s0_c23_n46_c;
                    stage1_col24[3] <= fa_s0_c23_n47_c;
                    stage1_col24[4] <= fa_s0_c24_n48_s;
                    stage1_col24[5] <= fa_s0_c24_n49_s;
                    stage1_col24[6] <= fa_s0_c24_n50_s;
                    stage1_col24[7] <= fa_s0_c24_n51_s;
                    stage1_col24[8] <= stage0_col24[12];
                    stage1_col24[9] <= stage0_col24[13];
                    stage1_col25[0] <= fa_s0_c24_n48_c;
                    stage1_col25[1] <= fa_s0_c24_n49_c;
                    stage1_col25[2] <= fa_s0_c24_n50_c;
                    stage1_col25[3] <= fa_s0_c24_n51_c;
                    stage1_col25[4] <= fa_s0_c25_n52_s;
                    stage1_col25[5] <= fa_s0_c25_n53_s;
                    stage1_col25[6] <= fa_s0_c25_n54_s;
                    stage1_col25[7] <= fa_s0_c25_n55_s;
                    stage1_col25[8] <= stage0_col25[12];
                    stage1_col26[0] <= fa_s0_c25_n52_c;
                    stage1_col26[1] <= fa_s0_c25_n53_c;
                    stage1_col26[2] <= fa_s0_c25_n54_c;
                    stage1_col26[3] <= fa_s0_c25_n55_c;
                    stage1_col26[4] <= fa_s0_c26_n56_s;
                    stage1_col26[5] <= fa_s0_c26_n57_s;
                    stage1_col26[6] <= fa_s0_c26_n58_s;
                    stage1_col26[7] <= fa_s0_c26_n59_s;
                    stage1_col26[8] <= fa_s0_c26_n60_s;
                    stage1_col27[0] <= fa_s0_c26_n56_c;
                    stage1_col27[1] <= fa_s0_c26_n57_c;
                    stage1_col27[2] <= fa_s0_c26_n58_c;
                    stage1_col27[3] <= fa_s0_c26_n59_c;
                    stage1_col27[4] <= fa_s0_c26_n60_c;
                    stage1_col27[5] <= fa_s0_c27_n61_s;
                    stage1_col27[6] <= fa_s0_c27_n62_s;
                    stage1_col27[7] <= fa_s0_c27_n63_s;
                    stage1_col27[8] <= fa_s0_c27_n64_s;
                    stage1_col27[9] <= stage0_col27[12];
                    stage1_col27[10] <= stage0_col27[13];
                    stage1_col28[0] <= fa_s0_c27_n61_c;
                    stage1_col28[1] <= fa_s0_c27_n62_c;
                    stage1_col28[2] <= fa_s0_c27_n63_c;
                    stage1_col28[3] <= fa_s0_c27_n64_c;
                    stage1_col28[4] <= fa_s0_c28_n65_s;
                    stage1_col28[5] <= fa_s0_c28_n66_s;
                    stage1_col28[6] <= fa_s0_c28_n67_s;
                    stage1_col28[7] <= fa_s0_c28_n68_s;
                    stage1_col28[8] <= fa_s0_c28_n69_s;
                    stage1_col28[9] <= stage0_col28[15];
                    stage1_col29[0] <= fa_s0_c28_n65_c;
                    stage1_col29[1] <= fa_s0_c28_n66_c;
                    stage1_col29[2] <= fa_s0_c28_n67_c;
                    stage1_col29[3] <= fa_s0_c28_n68_c;
                    stage1_col29[4] <= fa_s0_c28_n69_c;
                    stage1_col29[5] <= fa_s0_c29_n70_s;
                    stage1_col29[6] <= fa_s0_c29_n71_s;
                    stage1_col29[7] <= fa_s0_c29_n72_s;
                    stage1_col29[8] <= fa_s0_c29_n73_s;
                    stage1_col29[9] <= fa_s0_c29_n74_s;
                    stage1_col30[0] <= fa_s0_c29_n70_c;
                    stage1_col30[1] <= fa_s0_c29_n71_c;
                    stage1_col30[2] <= fa_s0_c29_n72_c;
                    stage1_col30[3] <= fa_s0_c29_n73_c;
                    stage1_col30[4] <= fa_s0_c29_n74_c;
                    stage1_col30[5] <= fa_s0_c30_n75_s;
                    stage1_col30[6] <= fa_s0_c30_n76_s;
                    stage1_col30[7] <= fa_s0_c30_n77_s;
                    stage1_col30[8] <= fa_s0_c30_n78_s;
                    stage1_col30[9] <= fa_s0_c30_n79_s;
                    stage1_col30[10] <= stage0_col30[15];
                    stage1_col30[11] <= stage0_col30[16];
                    stage1_col31[0] <= fa_s0_c30_n75_c;
                    stage1_col31[1] <= fa_s0_c30_n76_c;
                    stage1_col31[2] <= fa_s0_c30_n77_c;
                    stage1_col31[3] <= fa_s0_c30_n78_c;
                    stage1_col31[4] <= fa_s0_c30_n79_c;
                    stage1_col31[5] <= fa_s0_c31_n80_s;
                    stage1_col31[6] <= fa_s0_c31_n81_s;
                    stage1_col31[7] <= fa_s0_c31_n82_s;
                    stage1_col31[8] <= fa_s0_c31_n83_s;
                    stage1_col31[9] <= fa_s0_c31_n84_s;
                    stage1_col31[10] <= stage0_col31[15];
                    stage1_col32[0] <= fa_s0_c31_n80_c;
                    stage1_col32[1] <= fa_s0_c31_n81_c;
                    stage1_col32[2] <= fa_s0_c31_n82_c;
                    stage1_col32[3] <= fa_s0_c31_n83_c;
                    stage1_col32[4] <= fa_s0_c31_n84_c;
                    stage1_col32[5] <= fa_s0_c32_n85_s;
                    stage1_col32[6] <= fa_s0_c32_n86_s;
                    stage1_col32[7] <= fa_s0_c32_n87_s;
                    stage1_col32[8] <= fa_s0_c32_n88_s;
                    stage1_col32[9] <= fa_s0_c32_n89_s;
                    stage1_col32[10] <= fa_s0_c32_n90_s;
                    stage1_col33[0] <= fa_s0_c32_n85_c;
                    stage1_col33[1] <= fa_s0_c32_n86_c;
                    stage1_col33[2] <= fa_s0_c32_n87_c;
                    stage1_col33[3] <= fa_s0_c32_n88_c;
                    stage1_col33[4] <= fa_s0_c32_n89_c;
                    stage1_col33[5] <= fa_s0_c32_n90_c;
                    stage1_col33[6] <= fa_s0_c33_n91_s;
                    stage1_col33[7] <= fa_s0_c33_n92_s;
                    stage1_col33[8] <= fa_s0_c33_n93_s;
                    stage1_col33[9] <= fa_s0_c33_n94_s;
                    stage1_col33[10] <= fa_s0_c33_n95_s;
                    stage1_col33[11] <= stage0_col33[15];
                    stage1_col33[12] <= stage0_col33[16];
                    stage1_col34[0] <= fa_s0_c33_n91_c;
                    stage1_col34[1] <= fa_s0_c33_n92_c;
                    stage1_col34[2] <= fa_s0_c33_n93_c;
                    stage1_col34[3] <= fa_s0_c33_n94_c;
                    stage1_col34[4] <= fa_s0_c33_n95_c;
                    stage1_col34[5] <= fa_s0_c34_n96_s;
                    stage1_col34[6] <= fa_s0_c34_n97_s;
                    stage1_col34[7] <= fa_s0_c34_n98_s;
                    stage1_col34[8] <= fa_s0_c34_n99_s;
                    stage1_col34[9] <= fa_s0_c34_n100_s;
                    stage1_col34[10] <= fa_s0_c34_n101_s;
                    stage1_col34[11] <= stage0_col34[18];
                    stage1_col35[0] <= fa_s0_c34_n96_c;
                    stage1_col35[1] <= fa_s0_c34_n97_c;
                    stage1_col35[2] <= fa_s0_c34_n98_c;
                    stage1_col35[3] <= fa_s0_c34_n99_c;
                    stage1_col35[4] <= fa_s0_c34_n100_c;
                    stage1_col35[5] <= fa_s0_c34_n101_c;
                    stage1_col35[6] <= fa_s0_c35_n102_s;
                    stage1_col35[7] <= fa_s0_c35_n103_s;
                    stage1_col35[8] <= fa_s0_c35_n104_s;
                    stage1_col35[9] <= fa_s0_c35_n105_s;
                    stage1_col35[10] <= fa_s0_c35_n106_s;
                    stage1_col35[11] <= fa_s0_c35_n107_s;
                    stage1_col36[0] <= fa_s0_c35_n102_c;
                    stage1_col36[1] <= fa_s0_c35_n103_c;
                    stage1_col36[2] <= fa_s0_c35_n104_c;
                    stage1_col36[3] <= fa_s0_c35_n105_c;
                    stage1_col36[4] <= fa_s0_c35_n106_c;
                    stage1_col36[5] <= fa_s0_c35_n107_c;
                    stage1_col36[6] <= fa_s0_c36_n108_s;
                    stage1_col36[7] <= fa_s0_c36_n109_s;
                    stage1_col36[8] <= fa_s0_c36_n110_s;
                    stage1_col36[9] <= fa_s0_c36_n111_s;
                    stage1_col36[10] <= fa_s0_c36_n112_s;
                    stage1_col36[11] <= fa_s0_c36_n113_s;
                    stage1_col36[12] <= stage0_col36[18];
                    stage1_col36[13] <= stage0_col36[19];
                    stage1_col37[0] <= fa_s0_c36_n108_c;
                    stage1_col37[1] <= fa_s0_c36_n109_c;
                    stage1_col37[2] <= fa_s0_c36_n110_c;
                    stage1_col37[3] <= fa_s0_c36_n111_c;
                    stage1_col37[4] <= fa_s0_c36_n112_c;
                    stage1_col37[5] <= fa_s0_c36_n113_c;
                    stage1_col37[6] <= fa_s0_c37_n114_s;
                    stage1_col37[7] <= fa_s0_c37_n115_s;
                    stage1_col37[8] <= fa_s0_c37_n116_s;
                    stage1_col37[9] <= fa_s0_c37_n117_s;
                    stage1_col37[10] <= fa_s0_c37_n118_s;
                    stage1_col37[11] <= fa_s0_c37_n119_s;
                    stage1_col37[12] <= stage0_col37[18];
                    stage1_col38[0] <= fa_s0_c37_n114_c;
                    stage1_col38[1] <= fa_s0_c37_n115_c;
                    stage1_col38[2] <= fa_s0_c37_n116_c;
                    stage1_col38[3] <= fa_s0_c37_n117_c;
                    stage1_col38[4] <= fa_s0_c37_n118_c;
                    stage1_col38[5] <= fa_s0_c37_n119_c;
                    stage1_col38[6] <= fa_s0_c38_n120_s;
                    stage1_col38[7] <= fa_s0_c38_n121_s;
                    stage1_col38[8] <= fa_s0_c38_n122_s;
                    stage1_col38[9] <= fa_s0_c38_n123_s;
                    stage1_col38[10] <= fa_s0_c38_n124_s;
                    stage1_col38[11] <= fa_s0_c38_n125_s;
                    stage1_col38[12] <= fa_s0_c38_n126_s;
                    stage1_col39[0] <= fa_s0_c38_n120_c;
                    stage1_col39[1] <= fa_s0_c38_n121_c;
                    stage1_col39[2] <= fa_s0_c38_n122_c;
                    stage1_col39[3] <= fa_s0_c38_n123_c;
                    stage1_col39[4] <= fa_s0_c38_n124_c;
                    stage1_col39[5] <= fa_s0_c38_n125_c;
                    stage1_col39[6] <= fa_s0_c38_n126_c;
                    stage1_col39[7] <= fa_s0_c39_n127_s;
                    stage1_col39[8] <= fa_s0_c39_n128_s;
                    stage1_col39[9] <= fa_s0_c39_n129_s;
                    stage1_col39[10] <= fa_s0_c39_n130_s;
                    stage1_col39[11] <= fa_s0_c39_n131_s;
                    stage1_col39[12] <= fa_s0_c39_n132_s;
                    stage1_col39[13] <= stage0_col39[18];
                    stage1_col39[14] <= stage0_col39[19];
                    stage1_col40[0] <= fa_s0_c39_n127_c;
                    stage1_col40[1] <= fa_s0_c39_n128_c;
                    stage1_col40[2] <= fa_s0_c39_n129_c;
                    stage1_col40[3] <= fa_s0_c39_n130_c;
                    stage1_col40[4] <= fa_s0_c39_n131_c;
                    stage1_col40[5] <= fa_s0_c39_n132_c;
                    stage1_col40[6] <= fa_s0_c40_n133_s;
                    stage1_col40[7] <= fa_s0_c40_n134_s;
                    stage1_col40[8] <= fa_s0_c40_n135_s;
                    stage1_col40[9] <= fa_s0_c40_n136_s;
                    stage1_col40[10] <= fa_s0_c40_n137_s;
                    stage1_col40[11] <= fa_s0_c40_n138_s;
                    stage1_col40[12] <= fa_s0_c40_n139_s;
                    stage1_col40[13] <= stage0_col40[21];
                    stage1_col41[0] <= fa_s0_c40_n133_c;
                    stage1_col41[1] <= fa_s0_c40_n134_c;
                    stage1_col41[2] <= fa_s0_c40_n135_c;
                    stage1_col41[3] <= fa_s0_c40_n136_c;
                    stage1_col41[4] <= fa_s0_c40_n137_c;
                    stage1_col41[5] <= fa_s0_c40_n138_c;
                    stage1_col41[6] <= fa_s0_c40_n139_c;
                    stage1_col41[7] <= fa_s0_c41_n140_s;
                    stage1_col41[8] <= fa_s0_c41_n141_s;
                    stage1_col41[9] <= fa_s0_c41_n142_s;
                    stage1_col41[10] <= fa_s0_c41_n143_s;
                    stage1_col41[11] <= fa_s0_c41_n144_s;
                    stage1_col41[12] <= fa_s0_c41_n145_s;
                    stage1_col41[13] <= fa_s0_c41_n146_s;
                    stage1_col42[0] <= fa_s0_c41_n140_c;
                    stage1_col42[1] <= fa_s0_c41_n141_c;
                    stage1_col42[2] <= fa_s0_c41_n142_c;
                    stage1_col42[3] <= fa_s0_c41_n143_c;
                    stage1_col42[4] <= fa_s0_c41_n144_c;
                    stage1_col42[5] <= fa_s0_c41_n145_c;
                    stage1_col42[6] <= fa_s0_c41_n146_c;
                    stage1_col42[7] <= fa_s0_c42_n147_s;
                    stage1_col42[8] <= fa_s0_c42_n148_s;
                    stage1_col42[9] <= fa_s0_c42_n149_s;
                    stage1_col42[10] <= fa_s0_c42_n150_s;
                    stage1_col42[11] <= fa_s0_c42_n151_s;
                    stage1_col42[12] <= fa_s0_c42_n152_s;
                    stage1_col42[13] <= fa_s0_c42_n153_s;
                    stage1_col42[14] <= stage0_col42[21];
                    stage1_col42[15] <= stage0_col42[22];
                    stage1_col43[0] <= fa_s0_c42_n147_c;
                    stage1_col43[1] <= fa_s0_c42_n148_c;
                    stage1_col43[2] <= fa_s0_c42_n149_c;
                    stage1_col43[3] <= fa_s0_c42_n150_c;
                    stage1_col43[4] <= fa_s0_c42_n151_c;
                    stage1_col43[5] <= fa_s0_c42_n152_c;
                    stage1_col43[6] <= fa_s0_c42_n153_c;
                    stage1_col43[7] <= fa_s0_c43_n154_s;
                    stage1_col43[8] <= fa_s0_c43_n155_s;
                    stage1_col43[9] <= fa_s0_c43_n156_s;
                    stage1_col43[10] <= fa_s0_c43_n157_s;
                    stage1_col43[11] <= fa_s0_c43_n158_s;
                    stage1_col43[12] <= fa_s0_c43_n159_s;
                    stage1_col43[13] <= fa_s0_c43_n160_s;
                    stage1_col43[14] <= stage0_col43[21];
                    stage1_col44[0] <= fa_s0_c43_n154_c;
                    stage1_col44[1] <= fa_s0_c43_n155_c;
                    stage1_col44[2] <= fa_s0_c43_n156_c;
                    stage1_col44[3] <= fa_s0_c43_n157_c;
                    stage1_col44[4] <= fa_s0_c43_n158_c;
                    stage1_col44[5] <= fa_s0_c43_n159_c;
                    stage1_col44[6] <= fa_s0_c43_n160_c;
                    stage1_col44[7] <= fa_s0_c44_n161_s;
                    stage1_col44[8] <= fa_s0_c44_n162_s;
                    stage1_col44[9] <= fa_s0_c44_n163_s;
                    stage1_col44[10] <= fa_s0_c44_n164_s;
                    stage1_col44[11] <= fa_s0_c44_n165_s;
                    stage1_col44[12] <= fa_s0_c44_n166_s;
                    stage1_col44[13] <= fa_s0_c44_n167_s;
                    stage1_col44[14] <= fa_s0_c44_n168_s;
                    stage1_col45[0] <= fa_s0_c44_n161_c;
                    stage1_col45[1] <= fa_s0_c44_n162_c;
                    stage1_col45[2] <= fa_s0_c44_n163_c;
                    stage1_col45[3] <= fa_s0_c44_n164_c;
                    stage1_col45[4] <= fa_s0_c44_n165_c;
                    stage1_col45[5] <= fa_s0_c44_n166_c;
                    stage1_col45[6] <= fa_s0_c44_n167_c;
                    stage1_col45[7] <= fa_s0_c44_n168_c;
                    stage1_col45[8] <= fa_s0_c45_n169_s;
                    stage1_col45[9] <= fa_s0_c45_n170_s;
                    stage1_col45[10] <= fa_s0_c45_n171_s;
                    stage1_col45[11] <= fa_s0_c45_n172_s;
                    stage1_col45[12] <= fa_s0_c45_n173_s;
                    stage1_col45[13] <= fa_s0_c45_n174_s;
                    stage1_col45[14] <= fa_s0_c45_n175_s;
                    stage1_col45[15] <= stage0_col45[21];
                    stage1_col45[16] <= stage0_col45[22];
                    stage1_col46[0] <= fa_s0_c45_n169_c;
                    stage1_col46[1] <= fa_s0_c45_n170_c;
                    stage1_col46[2] <= fa_s0_c45_n171_c;
                    stage1_col46[3] <= fa_s0_c45_n172_c;
                    stage1_col46[4] <= fa_s0_c45_n173_c;
                    stage1_col46[5] <= fa_s0_c45_n174_c;
                    stage1_col46[6] <= fa_s0_c45_n175_c;
                    stage1_col46[7] <= fa_s0_c46_n176_s;
                    stage1_col46[8] <= fa_s0_c46_n177_s;
                    stage1_col46[9] <= fa_s0_c46_n178_s;
                    stage1_col46[10] <= fa_s0_c46_n179_s;
                    stage1_col46[11] <= fa_s0_c46_n180_s;
                    stage1_col46[12] <= fa_s0_c46_n181_s;
                    stage1_col46[13] <= fa_s0_c46_n182_s;
                    stage1_col46[14] <= fa_s0_c46_n183_s;
                    stage1_col46[15] <= stage0_col46[24];
                    stage1_col47[0] <= fa_s0_c46_n176_c;
                    stage1_col47[1] <= fa_s0_c46_n177_c;
                    stage1_col47[2] <= fa_s0_c46_n178_c;
                    stage1_col47[3] <= fa_s0_c46_n179_c;
                    stage1_col47[4] <= fa_s0_c46_n180_c;
                    stage1_col47[5] <= fa_s0_c46_n181_c;
                    stage1_col47[6] <= fa_s0_c46_n182_c;
                    stage1_col47[7] <= fa_s0_c46_n183_c;
                    stage1_col47[8] <= fa_s0_c47_n184_s;
                    stage1_col47[9] <= fa_s0_c47_n185_s;
                    stage1_col47[10] <= fa_s0_c47_n186_s;
                    stage1_col47[11] <= fa_s0_c47_n187_s;
                    stage1_col47[12] <= fa_s0_c47_n188_s;
                    stage1_col47[13] <= fa_s0_c47_n189_s;
                    stage1_col47[14] <= fa_s0_c47_n190_s;
                    stage1_col47[15] <= fa_s0_c47_n191_s;
                    stage1_col48[0] <= fa_s0_c47_n184_c;
                    stage1_col48[1] <= fa_s0_c47_n185_c;
                    stage1_col48[2] <= fa_s0_c47_n186_c;
                    stage1_col48[3] <= fa_s0_c47_n187_c;
                    stage1_col48[4] <= fa_s0_c47_n188_c;
                    stage1_col48[5] <= fa_s0_c47_n189_c;
                    stage1_col48[6] <= fa_s0_c47_n190_c;
                    stage1_col48[7] <= fa_s0_c47_n191_c;
                    stage1_col48[8] <= fa_s0_c48_n192_s;
                    stage1_col48[9] <= fa_s0_c48_n193_s;
                    stage1_col48[10] <= fa_s0_c48_n194_s;
                    stage1_col48[11] <= fa_s0_c48_n195_s;
                    stage1_col48[12] <= fa_s0_c48_n196_s;
                    stage1_col48[13] <= fa_s0_c48_n197_s;
                    stage1_col48[14] <= fa_s0_c48_n198_s;
                    stage1_col48[15] <= fa_s0_c48_n199_s;
                    stage1_col48[16] <= stage0_col48[24];
                    stage1_col48[17] <= stage0_col48[25];
                    stage1_col49[0] <= fa_s0_c48_n192_c;
                    stage1_col49[1] <= fa_s0_c48_n193_c;
                    stage1_col49[2] <= fa_s0_c48_n194_c;
                    stage1_col49[3] <= fa_s0_c48_n195_c;
                    stage1_col49[4] <= fa_s0_c48_n196_c;
                    stage1_col49[5] <= fa_s0_c48_n197_c;
                    stage1_col49[6] <= fa_s0_c48_n198_c;
                    stage1_col49[7] <= fa_s0_c48_n199_c;
                    stage1_col49[8] <= fa_s0_c49_n200_s;
                    stage1_col49[9] <= fa_s0_c49_n201_s;
                    stage1_col49[10] <= fa_s0_c49_n202_s;
                    stage1_col49[11] <= fa_s0_c49_n203_s;
                    stage1_col49[12] <= fa_s0_c49_n204_s;
                    stage1_col49[13] <= fa_s0_c49_n205_s;
                    stage1_col49[14] <= fa_s0_c49_n206_s;
                    stage1_col49[15] <= fa_s0_c49_n207_s;
                    stage1_col49[16] <= stage0_col49[24];
                    stage1_col50[0] <= fa_s0_c49_n200_c;
                    stage1_col50[1] <= fa_s0_c49_n201_c;
                    stage1_col50[2] <= fa_s0_c49_n202_c;
                    stage1_col50[3] <= fa_s0_c49_n203_c;
                    stage1_col50[4] <= fa_s0_c49_n204_c;
                    stage1_col50[5] <= fa_s0_c49_n205_c;
                    stage1_col50[6] <= fa_s0_c49_n206_c;
                    stage1_col50[7] <= fa_s0_c49_n207_c;
                    stage1_col50[8] <= fa_s0_c50_n208_s;
                    stage1_col50[9] <= fa_s0_c50_n209_s;
                    stage1_col50[10] <= fa_s0_c50_n210_s;
                    stage1_col50[11] <= fa_s0_c50_n211_s;
                    stage1_col50[12] <= fa_s0_c50_n212_s;
                    stage1_col50[13] <= fa_s0_c50_n213_s;
                    stage1_col50[14] <= fa_s0_c50_n214_s;
                    stage1_col50[15] <= fa_s0_c50_n215_s;
                    stage1_col50[16] <= fa_s0_c50_n216_s;
                    stage1_col51[0] <= fa_s0_c50_n208_c;
                    stage1_col51[1] <= fa_s0_c50_n209_c;
                    stage1_col51[2] <= fa_s0_c50_n210_c;
                    stage1_col51[3] <= fa_s0_c50_n211_c;
                    stage1_col51[4] <= fa_s0_c50_n212_c;
                    stage1_col51[5] <= fa_s0_c50_n213_c;
                    stage1_col51[6] <= fa_s0_c50_n214_c;
                    stage1_col51[7] <= fa_s0_c50_n215_c;
                    stage1_col51[8] <= fa_s0_c50_n216_c;
                    stage1_col51[9] <= fa_s0_c51_n217_s;
                    stage1_col51[10] <= fa_s0_c51_n218_s;
                    stage1_col51[11] <= fa_s0_c51_n219_s;
                    stage1_col51[12] <= fa_s0_c51_n220_s;
                    stage1_col51[13] <= fa_s0_c51_n221_s;
                    stage1_col51[14] <= fa_s0_c51_n222_s;
                    stage1_col51[15] <= fa_s0_c51_n223_s;
                    stage1_col51[16] <= fa_s0_c51_n224_s;
                    stage1_col51[17] <= stage0_col51[24];
                    stage1_col51[18] <= stage0_col51[25];
                    stage1_col52[0] <= fa_s0_c51_n217_c;
                    stage1_col52[1] <= fa_s0_c51_n218_c;
                    stage1_col52[2] <= fa_s0_c51_n219_c;
                    stage1_col52[3] <= fa_s0_c51_n220_c;
                    stage1_col52[4] <= fa_s0_c51_n221_c;
                    stage1_col52[5] <= fa_s0_c51_n222_c;
                    stage1_col52[6] <= fa_s0_c51_n223_c;
                    stage1_col52[7] <= fa_s0_c51_n224_c;
                    stage1_col52[8] <= fa_s0_c52_n225_s;
                    stage1_col52[9] <= fa_s0_c52_n226_s;
                    stage1_col52[10] <= fa_s0_c52_n227_s;
                    stage1_col52[11] <= fa_s0_c52_n228_s;
                    stage1_col52[12] <= fa_s0_c52_n229_s;
                    stage1_col52[13] <= fa_s0_c52_n230_s;
                    stage1_col52[14] <= fa_s0_c52_n231_s;
                    stage1_col52[15] <= fa_s0_c52_n232_s;
                    stage1_col52[16] <= fa_s0_c52_n233_s;
                    stage1_col52[17] <= stage0_col52[27];
                    stage1_col53[0] <= fa_s0_c52_n225_c;
                    stage1_col53[1] <= fa_s0_c52_n226_c;
                    stage1_col53[2] <= fa_s0_c52_n227_c;
                    stage1_col53[3] <= fa_s0_c52_n228_c;
                    stage1_col53[4] <= fa_s0_c52_n229_c;
                    stage1_col53[5] <= fa_s0_c52_n230_c;
                    stage1_col53[6] <= fa_s0_c52_n231_c;
                    stage1_col53[7] <= fa_s0_c52_n232_c;
                    stage1_col53[8] <= fa_s0_c52_n233_c;
                    stage1_col53[9] <= fa_s0_c53_n234_s;
                    stage1_col53[10] <= fa_s0_c53_n235_s;
                    stage1_col53[11] <= fa_s0_c53_n236_s;
                    stage1_col53[12] <= fa_s0_c53_n237_s;
                    stage1_col53[13] <= fa_s0_c53_n238_s;
                    stage1_col53[14] <= fa_s0_c53_n239_s;
                    stage1_col53[15] <= fa_s0_c53_n240_s;
                    stage1_col53[16] <= fa_s0_c53_n241_s;
                    stage1_col53[17] <= fa_s0_c53_n242_s;
                    stage1_col54[0] <= fa_s0_c53_n234_c;
                    stage1_col54[1] <= fa_s0_c53_n235_c;
                    stage1_col54[2] <= fa_s0_c53_n236_c;
                    stage1_col54[3] <= fa_s0_c53_n237_c;
                    stage1_col54[4] <= fa_s0_c53_n238_c;
                    stage1_col54[5] <= fa_s0_c53_n239_c;
                    stage1_col54[6] <= fa_s0_c53_n240_c;
                    stage1_col54[7] <= fa_s0_c53_n241_c;
                    stage1_col54[8] <= fa_s0_c53_n242_c;
                    stage1_col54[9] <= fa_s0_c54_n243_s;
                    stage1_col54[10] <= fa_s0_c54_n244_s;
                    stage1_col54[11] <= fa_s0_c54_n245_s;
                    stage1_col54[12] <= fa_s0_c54_n246_s;
                    stage1_col54[13] <= fa_s0_c54_n247_s;
                    stage1_col54[14] <= fa_s0_c54_n248_s;
                    stage1_col54[15] <= fa_s0_c54_n249_s;
                    stage1_col54[16] <= fa_s0_c54_n250_s;
                    stage1_col54[17] <= fa_s0_c54_n251_s;
                    stage1_col54[18] <= stage0_col54[27];
                    stage1_col54[19] <= stage0_col54[28];
                    stage1_col55[0] <= fa_s0_c54_n243_c;
                    stage1_col55[1] <= fa_s0_c54_n244_c;
                    stage1_col55[2] <= fa_s0_c54_n245_c;
                    stage1_col55[3] <= fa_s0_c54_n246_c;
                    stage1_col55[4] <= fa_s0_c54_n247_c;
                    stage1_col55[5] <= fa_s0_c54_n248_c;
                    stage1_col55[6] <= fa_s0_c54_n249_c;
                    stage1_col55[7] <= fa_s0_c54_n250_c;
                    stage1_col55[8] <= fa_s0_c54_n251_c;
                    stage1_col55[9] <= fa_s0_c55_n252_s;
                    stage1_col55[10] <= fa_s0_c55_n253_s;
                    stage1_col55[11] <= fa_s0_c55_n254_s;
                    stage1_col55[12] <= fa_s0_c55_n255_s;
                    stage1_col55[13] <= fa_s0_c55_n256_s;
                    stage1_col55[14] <= fa_s0_c55_n257_s;
                    stage1_col55[15] <= fa_s0_c55_n258_s;
                    stage1_col55[16] <= fa_s0_c55_n259_s;
                    stage1_col55[17] <= fa_s0_c55_n260_s;
                    stage1_col55[18] <= stage0_col55[27];
                    stage1_col56[0] <= fa_s0_c55_n252_c;
                    stage1_col56[1] <= fa_s0_c55_n253_c;
                    stage1_col56[2] <= fa_s0_c55_n254_c;
                    stage1_col56[3] <= fa_s0_c55_n255_c;
                    stage1_col56[4] <= fa_s0_c55_n256_c;
                    stage1_col56[5] <= fa_s0_c55_n257_c;
                    stage1_col56[6] <= fa_s0_c55_n258_c;
                    stage1_col56[7] <= fa_s0_c55_n259_c;
                    stage1_col56[8] <= fa_s0_c55_n260_c;
                    stage1_col56[9] <= fa_s0_c56_n261_s;
                    stage1_col56[10] <= fa_s0_c56_n262_s;
                    stage1_col56[11] <= fa_s0_c56_n263_s;
                    stage1_col56[12] <= fa_s0_c56_n264_s;
                    stage1_col56[13] <= fa_s0_c56_n265_s;
                    stage1_col56[14] <= fa_s0_c56_n266_s;
                    stage1_col56[15] <= fa_s0_c56_n267_s;
                    stage1_col56[16] <= fa_s0_c56_n268_s;
                    stage1_col56[17] <= fa_s0_c56_n269_s;
                    stage1_col56[18] <= fa_s0_c56_n270_s;
                    stage1_col57[0] <= fa_s0_c56_n261_c;
                    stage1_col57[1] <= fa_s0_c56_n262_c;
                    stage1_col57[2] <= fa_s0_c56_n263_c;
                    stage1_col57[3] <= fa_s0_c56_n264_c;
                    stage1_col57[4] <= fa_s0_c56_n265_c;
                    stage1_col57[5] <= fa_s0_c56_n266_c;
                    stage1_col57[6] <= fa_s0_c56_n267_c;
                    stage1_col57[7] <= fa_s0_c56_n268_c;
                    stage1_col57[8] <= fa_s0_c56_n269_c;
                    stage1_col57[9] <= fa_s0_c56_n270_c;
                    stage1_col57[10] <= fa_s0_c57_n271_s;
                    stage1_col57[11] <= fa_s0_c57_n272_s;
                    stage1_col57[12] <= fa_s0_c57_n273_s;
                    stage1_col57[13] <= fa_s0_c57_n274_s;
                    stage1_col57[14] <= fa_s0_c57_n275_s;
                    stage1_col57[15] <= fa_s0_c57_n276_s;
                    stage1_col57[16] <= fa_s0_c57_n277_s;
                    stage1_col57[17] <= fa_s0_c57_n278_s;
                    stage1_col57[18] <= fa_s0_c57_n279_s;
                    stage1_col57[19] <= stage0_col57[27];
                    stage1_col57[20] <= stage0_col57[28];
                    stage1_col58[0] <= fa_s0_c57_n271_c;
                    stage1_col58[1] <= fa_s0_c57_n272_c;
                    stage1_col58[2] <= fa_s0_c57_n273_c;
                    stage1_col58[3] <= fa_s0_c57_n274_c;
                    stage1_col58[4] <= fa_s0_c57_n275_c;
                    stage1_col58[5] <= fa_s0_c57_n276_c;
                    stage1_col58[6] <= fa_s0_c57_n277_c;
                    stage1_col58[7] <= fa_s0_c57_n278_c;
                    stage1_col58[8] <= fa_s0_c57_n279_c;
                    stage1_col58[9] <= fa_s0_c58_n280_s;
                    stage1_col58[10] <= fa_s0_c58_n281_s;
                    stage1_col58[11] <= fa_s0_c58_n282_s;
                    stage1_col58[12] <= fa_s0_c58_n283_s;
                    stage1_col58[13] <= fa_s0_c58_n284_s;
                    stage1_col58[14] <= fa_s0_c58_n285_s;
                    stage1_col58[15] <= fa_s0_c58_n286_s;
                    stage1_col58[16] <= fa_s0_c58_n287_s;
                    stage1_col58[17] <= fa_s0_c58_n288_s;
                    stage1_col58[18] <= fa_s0_c58_n289_s;
                    stage1_col58[19] <= stage0_col58[30];
                    stage1_col59[0] <= fa_s0_c58_n280_c;
                    stage1_col59[1] <= fa_s0_c58_n281_c;
                    stage1_col59[2] <= fa_s0_c58_n282_c;
                    stage1_col59[3] <= fa_s0_c58_n283_c;
                    stage1_col59[4] <= fa_s0_c58_n284_c;
                    stage1_col59[5] <= fa_s0_c58_n285_c;
                    stage1_col59[6] <= fa_s0_c58_n286_c;
                    stage1_col59[7] <= fa_s0_c58_n287_c;
                    stage1_col59[8] <= fa_s0_c58_n288_c;
                    stage1_col59[9] <= fa_s0_c58_n289_c;
                    stage1_col59[10] <= fa_s0_c59_n290_s;
                    stage1_col59[11] <= fa_s0_c59_n291_s;
                    stage1_col59[12] <= fa_s0_c59_n292_s;
                    stage1_col59[13] <= fa_s0_c59_n293_s;
                    stage1_col59[14] <= fa_s0_c59_n294_s;
                    stage1_col59[15] <= fa_s0_c59_n295_s;
                    stage1_col59[16] <= fa_s0_c59_n296_s;
                    stage1_col59[17] <= fa_s0_c59_n297_s;
                    stage1_col59[18] <= fa_s0_c59_n298_s;
                    stage1_col59[19] <= fa_s0_c59_n299_s;
                    stage1_col60[0] <= fa_s0_c59_n290_c;
                    stage1_col60[1] <= fa_s0_c59_n291_c;
                    stage1_col60[2] <= fa_s0_c59_n292_c;
                    stage1_col60[3] <= fa_s0_c59_n293_c;
                    stage1_col60[4] <= fa_s0_c59_n294_c;
                    stage1_col60[5] <= fa_s0_c59_n295_c;
                    stage1_col60[6] <= fa_s0_c59_n296_c;
                    stage1_col60[7] <= fa_s0_c59_n297_c;
                    stage1_col60[8] <= fa_s0_c59_n298_c;
                    stage1_col60[9] <= fa_s0_c59_n299_c;
                    stage1_col60[10] <= fa_s0_c60_n300_s;
                    stage1_col60[11] <= fa_s0_c60_n301_s;
                    stage1_col60[12] <= fa_s0_c60_n302_s;
                    stage1_col60[13] <= fa_s0_c60_n303_s;
                    stage1_col60[14] <= fa_s0_c60_n304_s;
                    stage1_col60[15] <= fa_s0_c60_n305_s;
                    stage1_col60[16] <= fa_s0_c60_n306_s;
                    stage1_col60[17] <= fa_s0_c60_n307_s;
                    stage1_col60[18] <= fa_s0_c60_n308_s;
                    stage1_col60[19] <= fa_s0_c60_n309_s;
                    stage1_col60[20] <= stage0_col60[30];
                    stage1_col60[21] <= stage0_col60[31];
                    stage1_col61[0] <= fa_s0_c60_n300_c;
                    stage1_col61[1] <= fa_s0_c60_n301_c;
                    stage1_col61[2] <= fa_s0_c60_n302_c;
                    stage1_col61[3] <= fa_s0_c60_n303_c;
                    stage1_col61[4] <= fa_s0_c60_n304_c;
                    stage1_col61[5] <= fa_s0_c60_n305_c;
                    stage1_col61[6] <= fa_s0_c60_n306_c;
                    stage1_col61[7] <= fa_s0_c60_n307_c;
                    stage1_col61[8] <= fa_s0_c60_n308_c;
                    stage1_col61[9] <= fa_s0_c60_n309_c;
                    stage1_col61[10] <= fa_s0_c61_n310_s;
                    stage1_col61[11] <= fa_s0_c61_n311_s;
                    stage1_col61[12] <= fa_s0_c61_n312_s;
                    stage1_col61[13] <= fa_s0_c61_n313_s;
                    stage1_col61[14] <= fa_s0_c61_n314_s;
                    stage1_col61[15] <= fa_s0_c61_n315_s;
                    stage1_col61[16] <= fa_s0_c61_n316_s;
                    stage1_col61[17] <= fa_s0_c61_n317_s;
                    stage1_col61[18] <= fa_s0_c61_n318_s;
                    stage1_col61[19] <= fa_s0_c61_n319_s;
                    stage1_col61[20] <= stage0_col61[30];
                    stage1_col62[0] <= fa_s0_c61_n310_c;
                    stage1_col62[1] <= fa_s0_c61_n311_c;
                    stage1_col62[2] <= fa_s0_c61_n312_c;
                    stage1_col62[3] <= fa_s0_c61_n313_c;
                    stage1_col62[4] <= fa_s0_c61_n314_c;
                    stage1_col62[5] <= fa_s0_c61_n315_c;
                    stage1_col62[6] <= fa_s0_c61_n316_c;
                    stage1_col62[7] <= fa_s0_c61_n317_c;
                    stage1_col62[8] <= fa_s0_c61_n318_c;
                    stage1_col62[9] <= fa_s0_c61_n319_c;
                    stage1_col62[10] <= fa_s0_c62_n320_s;
                    stage1_col62[11] <= fa_s0_c62_n321_s;
                    stage1_col62[12] <= fa_s0_c62_n322_s;
                    stage1_col62[13] <= fa_s0_c62_n323_s;
                    stage1_col62[14] <= fa_s0_c62_n324_s;
                    stage1_col62[15] <= fa_s0_c62_n325_s;
                    stage1_col62[16] <= fa_s0_c62_n326_s;
                    stage1_col62[17] <= fa_s0_c62_n327_s;
                    stage1_col62[18] <= fa_s0_c62_n328_s;
                    stage1_col62[19] <= fa_s0_c62_n329_s;
                    stage1_col62[20] <= fa_s0_c62_n330_s;
                    stage1_col63[0] <= fa_s0_c62_n320_c;
                    stage1_col63[1] <= fa_s0_c62_n321_c;
                    stage1_col63[2] <= fa_s0_c62_n322_c;
                    stage1_col63[3] <= fa_s0_c62_n323_c;
                    stage1_col63[4] <= fa_s0_c62_n324_c;
                    stage1_col63[5] <= fa_s0_c62_n325_c;
                    stage1_col63[6] <= fa_s0_c62_n326_c;
                    stage1_col63[7] <= fa_s0_c62_n327_c;
                    stage1_col63[8] <= fa_s0_c62_n328_c;
                    stage1_col63[9] <= fa_s0_c62_n329_c;
                    stage1_col63[10] <= fa_s0_c62_n330_c;
                    stage1_col63[11] <= fa_s0_c63_n331_s;
                    stage1_col63[12] <= fa_s0_c63_n332_s;
                    stage1_col63[13] <= fa_s0_c63_n333_s;
                    stage1_col63[14] <= fa_s0_c63_n334_s;
                    stage1_col63[15] <= fa_s0_c63_n335_s;
                    stage1_col63[16] <= fa_s0_c63_n336_s;
                    stage1_col63[17] <= fa_s0_c63_n337_s;
                    stage1_col63[18] <= fa_s0_c63_n338_s;
                    stage1_col63[19] <= fa_s0_c63_n339_s;
                    stage1_col63[20] <= fa_s0_c63_n340_s;
                    stage1_col63[21] <= stage0_col63[30];
                    stage1_col63[22] <= stage0_col63[31];
                    stage1_col64[0] <= fa_s0_c63_n331_c;
                    stage1_col64[1] <= fa_s0_c63_n332_c;
                    stage1_col64[2] <= fa_s0_c63_n333_c;
                    stage1_col64[3] <= fa_s0_c63_n334_c;
                    stage1_col64[4] <= fa_s0_c63_n335_c;
                    stage1_col64[5] <= fa_s0_c63_n336_c;
                    stage1_col64[6] <= fa_s0_c63_n337_c;
                    stage1_col64[7] <= fa_s0_c63_n338_c;
                    stage1_col64[8] <= fa_s0_c63_n339_c;
                    stage1_col64[9] <= fa_s0_c63_n340_c;
                    stage1_col64[10] <= fa_s0_c64_n341_s;
                    stage1_col64[11] <= fa_s0_c64_n342_s;
                    stage1_col64[12] <= fa_s0_c64_n343_s;
                    stage1_col64[13] <= fa_s0_c64_n344_s;
                    stage1_col64[14] <= fa_s0_c64_n345_s;
                    stage1_col64[15] <= fa_s0_c64_n346_s;
                    stage1_col64[16] <= fa_s0_c64_n347_s;
                    stage1_col64[17] <= fa_s0_c64_n348_s;
                    stage1_col64[18] <= fa_s0_c64_n349_s;
                    stage1_col64[19] <= fa_s0_c64_n350_s;
                    stage1_col64[20] <= fa_s0_c64_n351_s;
                    stage1_col65[0] <= fa_s0_c64_n341_c;
                    stage1_col65[1] <= fa_s0_c64_n342_c;
                    stage1_col65[2] <= fa_s0_c64_n343_c;
                    stage1_col65[3] <= fa_s0_c64_n344_c;
                    stage1_col65[4] <= fa_s0_c64_n345_c;
                    stage1_col65[5] <= fa_s0_c64_n346_c;
                    stage1_col65[6] <= fa_s0_c64_n347_c;
                    stage1_col65[7] <= fa_s0_c64_n348_c;
                    stage1_col65[8] <= fa_s0_c64_n349_c;
                    stage1_col65[9] <= fa_s0_c64_n350_c;
                    stage1_col65[10] <= fa_s0_c64_n351_c;
                    stage1_col65[11] <= fa_s0_c65_n352_s;
                    stage1_col65[12] <= fa_s0_c65_n353_s;
                    stage1_col65[13] <= fa_s0_c65_n354_s;
                    stage1_col65[14] <= fa_s0_c65_n355_s;
                    stage1_col65[15] <= fa_s0_c65_n356_s;
                    stage1_col65[16] <= fa_s0_c65_n357_s;
                    stage1_col65[17] <= fa_s0_c65_n358_s;
                    stage1_col65[18] <= fa_s0_c65_n359_s;
                    stage1_col65[19] <= fa_s0_c65_n360_s;
                    stage1_col65[20] <= fa_s0_c65_n361_s;
                    stage1_col65[21] <= stage0_col65[30];
                    stage1_col65[22] <= stage0_col65[31];
                    stage1_col66[0] <= fa_s0_c65_n352_c;
                    stage1_col66[1] <= fa_s0_c65_n353_c;
                    stage1_col66[2] <= fa_s0_c65_n354_c;
                    stage1_col66[3] <= fa_s0_c65_n355_c;
                    stage1_col66[4] <= fa_s0_c65_n356_c;
                    stage1_col66[5] <= fa_s0_c65_n357_c;
                    stage1_col66[6] <= fa_s0_c65_n358_c;
                    stage1_col66[7] <= fa_s0_c65_n359_c;
                    stage1_col66[8] <= fa_s0_c65_n360_c;
                    stage1_col66[9] <= fa_s0_c65_n361_c;
                    stage1_col66[10] <= fa_s0_c66_n362_s;
                    stage1_col66[11] <= fa_s0_c66_n363_s;
                    stage1_col66[12] <= fa_s0_c66_n364_s;
                    stage1_col66[13] <= fa_s0_c66_n365_s;
                    stage1_col66[14] <= fa_s0_c66_n366_s;
                    stage1_col66[15] <= fa_s0_c66_n367_s;
                    stage1_col66[16] <= fa_s0_c66_n368_s;
                    stage1_col66[17] <= fa_s0_c66_n369_s;
                    stage1_col66[18] <= fa_s0_c66_n370_s;
                    stage1_col66[19] <= fa_s0_c66_n371_s;
                    stage1_col66[20] <= fa_s0_c66_n372_s;
                    stage1_col67[0] <= fa_s0_c66_n362_c;
                    stage1_col67[1] <= fa_s0_c66_n363_c;
                    stage1_col67[2] <= fa_s0_c66_n364_c;
                    stage1_col67[3] <= fa_s0_c66_n365_c;
                    stage1_col67[4] <= fa_s0_c66_n366_c;
                    stage1_col67[5] <= fa_s0_c66_n367_c;
                    stage1_col67[6] <= fa_s0_c66_n368_c;
                    stage1_col67[7] <= fa_s0_c66_n369_c;
                    stage1_col67[8] <= fa_s0_c66_n370_c;
                    stage1_col67[9] <= fa_s0_c66_n371_c;
                    stage1_col67[10] <= fa_s0_c66_n372_c;
                    stage1_col67[11] <= fa_s0_c67_n373_s;
                    stage1_col67[12] <= fa_s0_c67_n374_s;
                    stage1_col67[13] <= fa_s0_c67_n375_s;
                    stage1_col67[14] <= fa_s0_c67_n376_s;
                    stage1_col67[15] <= fa_s0_c67_n377_s;
                    stage1_col67[16] <= fa_s0_c67_n378_s;
                    stage1_col67[17] <= fa_s0_c67_n379_s;
                    stage1_col67[18] <= fa_s0_c67_n380_s;
                    stage1_col67[19] <= fa_s0_c67_n381_s;
                    stage1_col67[20] <= fa_s0_c67_n382_s;
                    stage1_col67[21] <= stage0_col67[30];
                    stage1_col67[22] <= stage0_col67[31];
                    stage1_col68[0] <= fa_s0_c67_n373_c;
                    stage1_col68[1] <= fa_s0_c67_n374_c;
                    stage1_col68[2] <= fa_s0_c67_n375_c;
                    stage1_col68[3] <= fa_s0_c67_n376_c;
                    stage1_col68[4] <= fa_s0_c67_n377_c;
                    stage1_col68[5] <= fa_s0_c67_n378_c;
                    stage1_col68[6] <= fa_s0_c67_n379_c;
                    stage1_col68[7] <= fa_s0_c67_n380_c;
                    stage1_col68[8] <= fa_s0_c67_n381_c;
                    stage1_col68[9] <= fa_s0_c67_n382_c;
                    stage1_col68[10] <= fa_s0_c68_n383_s;
                    stage1_col68[11] <= fa_s0_c68_n384_s;
                    stage1_col68[12] <= fa_s0_c68_n385_s;
                    stage1_col68[13] <= fa_s0_c68_n386_s;
                    stage1_col68[14] <= fa_s0_c68_n387_s;
                    stage1_col68[15] <= fa_s0_c68_n388_s;
                    stage1_col68[16] <= fa_s0_c68_n389_s;
                    stage1_col68[17] <= fa_s0_c68_n390_s;
                    stage1_col68[18] <= fa_s0_c68_n391_s;
                    stage1_col68[19] <= fa_s0_c68_n392_s;
                    stage1_col68[20] <= fa_s0_c68_n393_s;
                    stage1_col69[0] <= fa_s0_c68_n383_c;
                    stage1_col69[1] <= fa_s0_c68_n384_c;
                    stage1_col69[2] <= fa_s0_c68_n385_c;
                    stage1_col69[3] <= fa_s0_c68_n386_c;
                    stage1_col69[4] <= fa_s0_c68_n387_c;
                    stage1_col69[5] <= fa_s0_c68_n388_c;
                    stage1_col69[6] <= fa_s0_c68_n389_c;
                    stage1_col69[7] <= fa_s0_c68_n390_c;
                    stage1_col69[8] <= fa_s0_c68_n391_c;
                    stage1_col69[9] <= fa_s0_c68_n392_c;
                    stage1_col69[10] <= fa_s0_c68_n393_c;
                    stage1_col69[11] <= fa_s0_c69_n394_s;
                    stage1_col69[12] <= fa_s0_c69_n395_s;
                    stage1_col69[13] <= fa_s0_c69_n396_s;
                    stage1_col69[14] <= fa_s0_c69_n397_s;
                    stage1_col69[15] <= fa_s0_c69_n398_s;
                    stage1_col69[16] <= fa_s0_c69_n399_s;
                    stage1_col69[17] <= fa_s0_c69_n400_s;
                    stage1_col69[18] <= fa_s0_c69_n401_s;
                    stage1_col69[19] <= fa_s0_c69_n402_s;
                    stage1_col69[20] <= fa_s0_c69_n403_s;
                    stage1_col69[21] <= stage0_col69[30];
                    stage1_col69[22] <= stage0_col69[31];
                    stage1_col70[0] <= fa_s0_c69_n394_c;
                    stage1_col70[1] <= fa_s0_c69_n395_c;
                    stage1_col70[2] <= fa_s0_c69_n396_c;
                    stage1_col70[3] <= fa_s0_c69_n397_c;
                    stage1_col70[4] <= fa_s0_c69_n398_c;
                    stage1_col70[5] <= fa_s0_c69_n399_c;
                    stage1_col70[6] <= fa_s0_c69_n400_c;
                    stage1_col70[7] <= fa_s0_c69_n401_c;
                    stage1_col70[8] <= fa_s0_c69_n402_c;
                    stage1_col70[9] <= fa_s0_c69_n403_c;
                    stage1_col70[10] <= fa_s0_c70_n404_s;
                    stage1_col70[11] <= fa_s0_c70_n405_s;
                    stage1_col70[12] <= fa_s0_c70_n406_s;
                    stage1_col70[13] <= fa_s0_c70_n407_s;
                    stage1_col70[14] <= fa_s0_c70_n408_s;
                    stage1_col70[15] <= fa_s0_c70_n409_s;
                    stage1_col70[16] <= fa_s0_c70_n410_s;
                    stage1_col70[17] <= fa_s0_c70_n411_s;
                    stage1_col70[18] <= fa_s0_c70_n412_s;
                    stage1_col70[19] <= fa_s0_c70_n413_s;
                    stage1_col70[20] <= fa_s0_c70_n414_s;
                    stage1_col71[0] <= fa_s0_c70_n404_c;
                    stage1_col71[1] <= fa_s0_c70_n405_c;
                    stage1_col71[2] <= fa_s0_c70_n406_c;
                    stage1_col71[3] <= fa_s0_c70_n407_c;
                    stage1_col71[4] <= fa_s0_c70_n408_c;
                    stage1_col71[5] <= fa_s0_c70_n409_c;
                    stage1_col71[6] <= fa_s0_c70_n410_c;
                    stage1_col71[7] <= fa_s0_c70_n411_c;
                    stage1_col71[8] <= fa_s0_c70_n412_c;
                    stage1_col71[9] <= fa_s0_c70_n413_c;
                    stage1_col71[10] <= fa_s0_c70_n414_c;
                    stage1_col71[11] <= fa_s0_c71_n415_s;
                    stage1_col71[12] <= fa_s0_c71_n416_s;
                    stage1_col71[13] <= fa_s0_c71_n417_s;
                    stage1_col71[14] <= fa_s0_c71_n418_s;
                    stage1_col71[15] <= fa_s0_c71_n419_s;
                    stage1_col71[16] <= fa_s0_c71_n420_s;
                    stage1_col71[17] <= fa_s0_c71_n421_s;
                    stage1_col71[18] <= fa_s0_c71_n422_s;
                    stage1_col71[19] <= fa_s0_c71_n423_s;
                    stage1_col71[20] <= fa_s0_c71_n424_s;
                    stage1_col71[21] <= stage0_col71[30];
                    stage1_col71[22] <= stage0_col71[31];
                    stage1_col72[0] <= fa_s0_c71_n415_c;
                    stage1_col72[1] <= fa_s0_c71_n416_c;
                    stage1_col72[2] <= fa_s0_c71_n417_c;
                    stage1_col72[3] <= fa_s0_c71_n418_c;
                    stage1_col72[4] <= fa_s0_c71_n419_c;
                    stage1_col72[5] <= fa_s0_c71_n420_c;
                    stage1_col72[6] <= fa_s0_c71_n421_c;
                    stage1_col72[7] <= fa_s0_c71_n422_c;
                    stage1_col72[8] <= fa_s0_c71_n423_c;
                    stage1_col72[9] <= fa_s0_c71_n424_c;
                    stage1_col72[10] <= fa_s0_c72_n425_s;
                    stage1_col72[11] <= fa_s0_c72_n426_s;
                    stage1_col72[12] <= fa_s0_c72_n427_s;
                    stage1_col72[13] <= fa_s0_c72_n428_s;
                    stage1_col72[14] <= fa_s0_c72_n429_s;
                    stage1_col72[15] <= fa_s0_c72_n430_s;
                    stage1_col72[16] <= fa_s0_c72_n431_s;
                    stage1_col72[17] <= fa_s0_c72_n432_s;
                    stage1_col72[18] <= fa_s0_c72_n433_s;
                    stage1_col72[19] <= fa_s0_c72_n434_s;
                    stage1_col72[20] <= fa_s0_c72_n435_s;
                    stage1_col73[0] <= fa_s0_c72_n425_c;
                    stage1_col73[1] <= fa_s0_c72_n426_c;
                    stage1_col73[2] <= fa_s0_c72_n427_c;
                    stage1_col73[3] <= fa_s0_c72_n428_c;
                    stage1_col73[4] <= fa_s0_c72_n429_c;
                    stage1_col73[5] <= fa_s0_c72_n430_c;
                    stage1_col73[6] <= fa_s0_c72_n431_c;
                    stage1_col73[7] <= fa_s0_c72_n432_c;
                    stage1_col73[8] <= fa_s0_c72_n433_c;
                    stage1_col73[9] <= fa_s0_c72_n434_c;
                    stage1_col73[10] <= fa_s0_c72_n435_c;
                    stage1_col73[11] <= fa_s0_c73_n436_s;
                    stage1_col73[12] <= fa_s0_c73_n437_s;
                    stage1_col73[13] <= fa_s0_c73_n438_s;
                    stage1_col73[14] <= fa_s0_c73_n439_s;
                    stage1_col73[15] <= fa_s0_c73_n440_s;
                    stage1_col73[16] <= fa_s0_c73_n441_s;
                    stage1_col73[17] <= fa_s0_c73_n442_s;
                    stage1_col73[18] <= fa_s0_c73_n443_s;
                    stage1_col73[19] <= fa_s0_c73_n444_s;
                    stage1_col73[20] <= fa_s0_c73_n445_s;
                    stage1_col73[21] <= stage0_col73[30];
                    stage1_col73[22] <= stage0_col73[31];
                    stage1_col74[0] <= fa_s0_c73_n436_c;
                    stage1_col74[1] <= fa_s0_c73_n437_c;
                    stage1_col74[2] <= fa_s0_c73_n438_c;
                    stage1_col74[3] <= fa_s0_c73_n439_c;
                    stage1_col74[4] <= fa_s0_c73_n440_c;
                    stage1_col74[5] <= fa_s0_c73_n441_c;
                    stage1_col74[6] <= fa_s0_c73_n442_c;
                    stage1_col74[7] <= fa_s0_c73_n443_c;
                    stage1_col74[8] <= fa_s0_c73_n444_c;
                    stage1_col74[9] <= fa_s0_c73_n445_c;
                    stage1_col74[10] <= fa_s0_c74_n446_s;
                    stage1_col74[11] <= fa_s0_c74_n447_s;
                    stage1_col74[12] <= fa_s0_c74_n448_s;
                    stage1_col74[13] <= fa_s0_c74_n449_s;
                    stage1_col74[14] <= fa_s0_c74_n450_s;
                    stage1_col74[15] <= fa_s0_c74_n451_s;
                    stage1_col74[16] <= fa_s0_c74_n452_s;
                    stage1_col74[17] <= fa_s0_c74_n453_s;
                    stage1_col74[18] <= fa_s0_c74_n454_s;
                    stage1_col74[19] <= fa_s0_c74_n455_s;
                    stage1_col74[20] <= fa_s0_c74_n456_s;
                    stage1_col75[0] <= fa_s0_c74_n446_c;
                    stage1_col75[1] <= fa_s0_c74_n447_c;
                    stage1_col75[2] <= fa_s0_c74_n448_c;
                    stage1_col75[3] <= fa_s0_c74_n449_c;
                    stage1_col75[4] <= fa_s0_c74_n450_c;
                    stage1_col75[5] <= fa_s0_c74_n451_c;
                    stage1_col75[6] <= fa_s0_c74_n452_c;
                    stage1_col75[7] <= fa_s0_c74_n453_c;
                    stage1_col75[8] <= fa_s0_c74_n454_c;
                    stage1_col75[9] <= fa_s0_c74_n455_c;
                    stage1_col75[10] <= fa_s0_c74_n456_c;
                    stage1_col75[11] <= fa_s0_c75_n457_s;
                    stage1_col75[12] <= fa_s0_c75_n458_s;
                    stage1_col75[13] <= fa_s0_c75_n459_s;
                    stage1_col75[14] <= fa_s0_c75_n460_s;
                    stage1_col75[15] <= fa_s0_c75_n461_s;
                    stage1_col75[16] <= fa_s0_c75_n462_s;
                    stage1_col75[17] <= fa_s0_c75_n463_s;
                    stage1_col75[18] <= fa_s0_c75_n464_s;
                    stage1_col75[19] <= fa_s0_c75_n465_s;
                    stage1_col75[20] <= fa_s0_c75_n466_s;
                    stage1_col75[21] <= stage0_col75[30];
                    stage1_col75[22] <= stage0_col75[31];
                    stage1_col76[0] <= fa_s0_c75_n457_c;
                    stage1_col76[1] <= fa_s0_c75_n458_c;
                    stage1_col76[2] <= fa_s0_c75_n459_c;
                    stage1_col76[3] <= fa_s0_c75_n460_c;
                    stage1_col76[4] <= fa_s0_c75_n461_c;
                    stage1_col76[5] <= fa_s0_c75_n462_c;
                    stage1_col76[6] <= fa_s0_c75_n463_c;
                    stage1_col76[7] <= fa_s0_c75_n464_c;
                    stage1_col76[8] <= fa_s0_c75_n465_c;
                    stage1_col76[9] <= fa_s0_c75_n466_c;
                    stage1_col76[10] <= fa_s0_c76_n467_s;
                    stage1_col76[11] <= fa_s0_c76_n468_s;
                    stage1_col76[12] <= fa_s0_c76_n469_s;
                    stage1_col76[13] <= fa_s0_c76_n470_s;
                    stage1_col76[14] <= fa_s0_c76_n471_s;
                    stage1_col76[15] <= fa_s0_c76_n472_s;
                    stage1_col76[16] <= fa_s0_c76_n473_s;
                    stage1_col76[17] <= fa_s0_c76_n474_s;
                    stage1_col76[18] <= fa_s0_c76_n475_s;
                    stage1_col76[19] <= fa_s0_c76_n476_s;
                    stage1_col76[20] <= fa_s0_c76_n477_s;
                    stage1_col77[0] <= fa_s0_c76_n467_c;
                    stage1_col77[1] <= fa_s0_c76_n468_c;
                    stage1_col77[2] <= fa_s0_c76_n469_c;
                    stage1_col77[3] <= fa_s0_c76_n470_c;
                    stage1_col77[4] <= fa_s0_c76_n471_c;
                    stage1_col77[5] <= fa_s0_c76_n472_c;
                    stage1_col77[6] <= fa_s0_c76_n473_c;
                    stage1_col77[7] <= fa_s0_c76_n474_c;
                    stage1_col77[8] <= fa_s0_c76_n475_c;
                    stage1_col77[9] <= fa_s0_c76_n476_c;
                    stage1_col77[10] <= fa_s0_c76_n477_c;
                    stage1_col77[11] <= fa_s0_c77_n478_s;
                    stage1_col77[12] <= fa_s0_c77_n479_s;
                    stage1_col77[13] <= fa_s0_c77_n480_s;
                    stage1_col77[14] <= fa_s0_c77_n481_s;
                    stage1_col77[15] <= fa_s0_c77_n482_s;
                    stage1_col77[16] <= fa_s0_c77_n483_s;
                    stage1_col77[17] <= fa_s0_c77_n484_s;
                    stage1_col77[18] <= fa_s0_c77_n485_s;
                    stage1_col77[19] <= fa_s0_c77_n486_s;
                    stage1_col77[20] <= fa_s0_c77_n487_s;
                    stage1_col77[21] <= stage0_col77[30];
                    stage1_col77[22] <= stage0_col77[31];
                    stage1_col78[0] <= fa_s0_c77_n478_c;
                    stage1_col78[1] <= fa_s0_c77_n479_c;
                    stage1_col78[2] <= fa_s0_c77_n480_c;
                    stage1_col78[3] <= fa_s0_c77_n481_c;
                    stage1_col78[4] <= fa_s0_c77_n482_c;
                    stage1_col78[5] <= fa_s0_c77_n483_c;
                    stage1_col78[6] <= fa_s0_c77_n484_c;
                    stage1_col78[7] <= fa_s0_c77_n485_c;
                    stage1_col78[8] <= fa_s0_c77_n486_c;
                    stage1_col78[9] <= fa_s0_c77_n487_c;
                    stage1_col78[10] <= fa_s0_c78_n488_s;
                    stage1_col78[11] <= fa_s0_c78_n489_s;
                    stage1_col78[12] <= fa_s0_c78_n490_s;
                    stage1_col78[13] <= fa_s0_c78_n491_s;
                    stage1_col78[14] <= fa_s0_c78_n492_s;
                    stage1_col78[15] <= fa_s0_c78_n493_s;
                    stage1_col78[16] <= fa_s0_c78_n494_s;
                    stage1_col78[17] <= fa_s0_c78_n495_s;
                    stage1_col78[18] <= fa_s0_c78_n496_s;
                    stage1_col78[19] <= fa_s0_c78_n497_s;
                    stage1_col78[20] <= fa_s0_c78_n498_s;
                    stage1_col79[0] <= fa_s0_c78_n488_c;
                    stage1_col79[1] <= fa_s0_c78_n489_c;
                    stage1_col79[2] <= fa_s0_c78_n490_c;
                    stage1_col79[3] <= fa_s0_c78_n491_c;
                    stage1_col79[4] <= fa_s0_c78_n492_c;
                    stage1_col79[5] <= fa_s0_c78_n493_c;
                    stage1_col79[6] <= fa_s0_c78_n494_c;
                    stage1_col79[7] <= fa_s0_c78_n495_c;
                    stage1_col79[8] <= fa_s0_c78_n496_c;
                    stage1_col79[9] <= fa_s0_c78_n497_c;
                    stage1_col79[10] <= fa_s0_c78_n498_c;
                    stage1_col79[11] <= fa_s0_c79_n499_s;
                    stage1_col79[12] <= fa_s0_c79_n500_s;
                    stage1_col79[13] <= fa_s0_c79_n501_s;
                    stage1_col79[14] <= fa_s0_c79_n502_s;
                    stage1_col79[15] <= fa_s0_c79_n503_s;
                    stage1_col79[16] <= fa_s0_c79_n504_s;
                    stage1_col79[17] <= fa_s0_c79_n505_s;
                    stage1_col79[18] <= fa_s0_c79_n506_s;
                    stage1_col79[19] <= fa_s0_c79_n507_s;
                    stage1_col79[20] <= fa_s0_c79_n508_s;
                    stage1_col79[21] <= stage0_col79[30];
                    stage1_col79[22] <= stage0_col79[31];
                    stage1_col80[0] <= fa_s0_c79_n499_c;
                    stage1_col80[1] <= fa_s0_c79_n500_c;
                    stage1_col80[2] <= fa_s0_c79_n501_c;
                    stage1_col80[3] <= fa_s0_c79_n502_c;
                    stage1_col80[4] <= fa_s0_c79_n503_c;
                    stage1_col80[5] <= fa_s0_c79_n504_c;
                    stage1_col80[6] <= fa_s0_c79_n505_c;
                    stage1_col80[7] <= fa_s0_c79_n506_c;
                    stage1_col80[8] <= fa_s0_c79_n507_c;
                    stage1_col80[9] <= fa_s0_c79_n508_c;
                    stage1_col80[10] <= fa_s0_c80_n509_s;
                    stage1_col80[11] <= fa_s0_c80_n510_s;
                    stage1_col80[12] <= fa_s0_c80_n511_s;
                    stage1_col80[13] <= fa_s0_c80_n512_s;
                    stage1_col80[14] <= fa_s0_c80_n513_s;
                    stage1_col80[15] <= fa_s0_c80_n514_s;
                    stage1_col80[16] <= fa_s0_c80_n515_s;
                    stage1_col80[17] <= fa_s0_c80_n516_s;
                    stage1_col80[18] <= fa_s0_c80_n517_s;
                    stage1_col80[19] <= fa_s0_c80_n518_s;
                    stage1_col80[20] <= fa_s0_c80_n519_s;
                    stage1_col81[0] <= fa_s0_c80_n509_c;
                    stage1_col81[1] <= fa_s0_c80_n510_c;
                    stage1_col81[2] <= fa_s0_c80_n511_c;
                    stage1_col81[3] <= fa_s0_c80_n512_c;
                    stage1_col81[4] <= fa_s0_c80_n513_c;
                    stage1_col81[5] <= fa_s0_c80_n514_c;
                    stage1_col81[6] <= fa_s0_c80_n515_c;
                    stage1_col81[7] <= fa_s0_c80_n516_c;
                    stage1_col81[8] <= fa_s0_c80_n517_c;
                    stage1_col81[9] <= fa_s0_c80_n518_c;
                    stage1_col81[10] <= fa_s0_c80_n519_c;
                    stage1_col81[11] <= fa_s0_c81_n520_s;
                    stage1_col81[12] <= fa_s0_c81_n521_s;
                    stage1_col81[13] <= fa_s0_c81_n522_s;
                    stage1_col81[14] <= fa_s0_c81_n523_s;
                    stage1_col81[15] <= fa_s0_c81_n524_s;
                    stage1_col81[16] <= fa_s0_c81_n525_s;
                    stage1_col81[17] <= fa_s0_c81_n526_s;
                    stage1_col81[18] <= fa_s0_c81_n527_s;
                    stage1_col81[19] <= fa_s0_c81_n528_s;
                    stage1_col81[20] <= fa_s0_c81_n529_s;
                    stage1_col81[21] <= stage0_col81[30];
                    stage1_col81[22] <= stage0_col81[31];
                    stage1_col82[0] <= fa_s0_c81_n520_c;
                    stage1_col82[1] <= fa_s0_c81_n521_c;
                    stage1_col82[2] <= fa_s0_c81_n522_c;
                    stage1_col82[3] <= fa_s0_c81_n523_c;
                    stage1_col82[4] <= fa_s0_c81_n524_c;
                    stage1_col82[5] <= fa_s0_c81_n525_c;
                    stage1_col82[6] <= fa_s0_c81_n526_c;
                    stage1_col82[7] <= fa_s0_c81_n527_c;
                    stage1_col82[8] <= fa_s0_c81_n528_c;
                    stage1_col82[9] <= fa_s0_c81_n529_c;
                    stage1_col82[10] <= fa_s0_c82_n530_s;
                    stage1_col82[11] <= fa_s0_c82_n531_s;
                    stage1_col82[12] <= fa_s0_c82_n532_s;
                    stage1_col82[13] <= fa_s0_c82_n533_s;
                    stage1_col82[14] <= fa_s0_c82_n534_s;
                    stage1_col82[15] <= fa_s0_c82_n535_s;
                    stage1_col82[16] <= fa_s0_c82_n536_s;
                    stage1_col82[17] <= fa_s0_c82_n537_s;
                    stage1_col82[18] <= fa_s0_c82_n538_s;
                    stage1_col82[19] <= fa_s0_c82_n539_s;
                    stage1_col82[20] <= fa_s0_c82_n540_s;
                    stage1_col83[0] <= fa_s0_c82_n530_c;
                    stage1_col83[1] <= fa_s0_c82_n531_c;
                    stage1_col83[2] <= fa_s0_c82_n532_c;
                    stage1_col83[3] <= fa_s0_c82_n533_c;
                    stage1_col83[4] <= fa_s0_c82_n534_c;
                    stage1_col83[5] <= fa_s0_c82_n535_c;
                    stage1_col83[6] <= fa_s0_c82_n536_c;
                    stage1_col83[7] <= fa_s0_c82_n537_c;
                    stage1_col83[8] <= fa_s0_c82_n538_c;
                    stage1_col83[9] <= fa_s0_c82_n539_c;
                    stage1_col83[10] <= fa_s0_c82_n540_c;
                    stage1_col83[11] <= fa_s0_c83_n541_s;
                    stage1_col83[12] <= fa_s0_c83_n542_s;
                    stage1_col83[13] <= fa_s0_c83_n543_s;
                    stage1_col83[14] <= fa_s0_c83_n544_s;
                    stage1_col83[15] <= fa_s0_c83_n545_s;
                    stage1_col83[16] <= fa_s0_c83_n546_s;
                    stage1_col83[17] <= fa_s0_c83_n547_s;
                    stage1_col83[18] <= fa_s0_c83_n548_s;
                    stage1_col83[19] <= fa_s0_c83_n549_s;
                    stage1_col83[20] <= fa_s0_c83_n550_s;
                    stage1_col83[21] <= stage0_col83[30];
                    stage1_col83[22] <= stage0_col83[31];
                    stage1_col84[0] <= fa_s0_c83_n541_c;
                    stage1_col84[1] <= fa_s0_c83_n542_c;
                    stage1_col84[2] <= fa_s0_c83_n543_c;
                    stage1_col84[3] <= fa_s0_c83_n544_c;
                    stage1_col84[4] <= fa_s0_c83_n545_c;
                    stage1_col84[5] <= fa_s0_c83_n546_c;
                    stage1_col84[6] <= fa_s0_c83_n547_c;
                    stage1_col84[7] <= fa_s0_c83_n548_c;
                    stage1_col84[8] <= fa_s0_c83_n549_c;
                    stage1_col84[9] <= fa_s0_c83_n550_c;
                    stage1_col84[10] <= fa_s0_c84_n551_s;
                    stage1_col84[11] <= fa_s0_c84_n552_s;
                    stage1_col84[12] <= fa_s0_c84_n553_s;
                    stage1_col84[13] <= fa_s0_c84_n554_s;
                    stage1_col84[14] <= fa_s0_c84_n555_s;
                    stage1_col84[15] <= fa_s0_c84_n556_s;
                    stage1_col84[16] <= fa_s0_c84_n557_s;
                    stage1_col84[17] <= fa_s0_c84_n558_s;
                    stage1_col84[18] <= fa_s0_c84_n559_s;
                    stage1_col84[19] <= fa_s0_c84_n560_s;
                    stage1_col84[20] <= fa_s0_c84_n561_s;
                    stage1_col85[0] <= fa_s0_c84_n551_c;
                    stage1_col85[1] <= fa_s0_c84_n552_c;
                    stage1_col85[2] <= fa_s0_c84_n553_c;
                    stage1_col85[3] <= fa_s0_c84_n554_c;
                    stage1_col85[4] <= fa_s0_c84_n555_c;
                    stage1_col85[5] <= fa_s0_c84_n556_c;
                    stage1_col85[6] <= fa_s0_c84_n557_c;
                    stage1_col85[7] <= fa_s0_c84_n558_c;
                    stage1_col85[8] <= fa_s0_c84_n559_c;
                    stage1_col85[9] <= fa_s0_c84_n560_c;
                    stage1_col85[10] <= fa_s0_c84_n561_c;
                    stage1_col85[11] <= fa_s0_c85_n562_s;
                    stage1_col85[12] <= fa_s0_c85_n563_s;
                    stage1_col85[13] <= fa_s0_c85_n564_s;
                    stage1_col85[14] <= fa_s0_c85_n565_s;
                    stage1_col85[15] <= fa_s0_c85_n566_s;
                    stage1_col85[16] <= fa_s0_c85_n567_s;
                    stage1_col85[17] <= fa_s0_c85_n568_s;
                    stage1_col85[18] <= fa_s0_c85_n569_s;
                    stage1_col85[19] <= fa_s0_c85_n570_s;
                    stage1_col85[20] <= fa_s0_c85_n571_s;
                    stage1_col85[21] <= stage0_col85[30];
                    stage1_col85[22] <= stage0_col85[31];
                    stage1_col86[0] <= fa_s0_c85_n562_c;
                    stage1_col86[1] <= fa_s0_c85_n563_c;
                    stage1_col86[2] <= fa_s0_c85_n564_c;
                    stage1_col86[3] <= fa_s0_c85_n565_c;
                    stage1_col86[4] <= fa_s0_c85_n566_c;
                    stage1_col86[5] <= fa_s0_c85_n567_c;
                    stage1_col86[6] <= fa_s0_c85_n568_c;
                    stage1_col86[7] <= fa_s0_c85_n569_c;
                    stage1_col86[8] <= fa_s0_c85_n570_c;
                    stage1_col86[9] <= fa_s0_c85_n571_c;
                    stage1_col86[10] <= fa_s0_c86_n572_s;
                    stage1_col86[11] <= fa_s0_c86_n573_s;
                    stage1_col86[12] <= fa_s0_c86_n574_s;
                    stage1_col86[13] <= fa_s0_c86_n575_s;
                    stage1_col86[14] <= fa_s0_c86_n576_s;
                    stage1_col86[15] <= fa_s0_c86_n577_s;
                    stage1_col86[16] <= fa_s0_c86_n578_s;
                    stage1_col86[17] <= fa_s0_c86_n579_s;
                    stage1_col86[18] <= fa_s0_c86_n580_s;
                    stage1_col86[19] <= fa_s0_c86_n581_s;
                    stage1_col86[20] <= fa_s0_c86_n582_s;
                    stage1_col87[0] <= fa_s0_c86_n572_c;
                    stage1_col87[1] <= fa_s0_c86_n573_c;
                    stage1_col87[2] <= fa_s0_c86_n574_c;
                    stage1_col87[3] <= fa_s0_c86_n575_c;
                    stage1_col87[4] <= fa_s0_c86_n576_c;
                    stage1_col87[5] <= fa_s0_c86_n577_c;
                    stage1_col87[6] <= fa_s0_c86_n578_c;
                    stage1_col87[7] <= fa_s0_c86_n579_c;
                    stage1_col87[8] <= fa_s0_c86_n580_c;
                    stage1_col87[9] <= fa_s0_c86_n581_c;
                    stage1_col87[10] <= fa_s0_c86_n582_c;
                    stage1_col87[11] <= fa_s0_c87_n583_s;
                    stage1_col87[12] <= fa_s0_c87_n584_s;
                    stage1_col87[13] <= fa_s0_c87_n585_s;
                    stage1_col87[14] <= fa_s0_c87_n586_s;
                    stage1_col87[15] <= fa_s0_c87_n587_s;
                    stage1_col87[16] <= fa_s0_c87_n588_s;
                    stage1_col87[17] <= fa_s0_c87_n589_s;
                    stage1_col87[18] <= fa_s0_c87_n590_s;
                    stage1_col87[19] <= fa_s0_c87_n591_s;
                    stage1_col87[20] <= fa_s0_c87_n592_s;
                    stage1_col87[21] <= stage0_col87[30];
                    stage1_col87[22] <= stage0_col87[31];
                    stage1_col88[0] <= fa_s0_c87_n583_c;
                    stage1_col88[1] <= fa_s0_c87_n584_c;
                    stage1_col88[2] <= fa_s0_c87_n585_c;
                    stage1_col88[3] <= fa_s0_c87_n586_c;
                    stage1_col88[4] <= fa_s0_c87_n587_c;
                    stage1_col88[5] <= fa_s0_c87_n588_c;
                    stage1_col88[6] <= fa_s0_c87_n589_c;
                    stage1_col88[7] <= fa_s0_c87_n590_c;
                    stage1_col88[8] <= fa_s0_c87_n591_c;
                    stage1_col88[9] <= fa_s0_c87_n592_c;
                    stage1_col88[10] <= fa_s0_c88_n593_s;
                    stage1_col88[11] <= fa_s0_c88_n594_s;
                    stage1_col88[12] <= fa_s0_c88_n595_s;
                    stage1_col88[13] <= fa_s0_c88_n596_s;
                    stage1_col88[14] <= fa_s0_c88_n597_s;
                    stage1_col88[15] <= fa_s0_c88_n598_s;
                    stage1_col88[16] <= fa_s0_c88_n599_s;
                    stage1_col88[17] <= fa_s0_c88_n600_s;
                    stage1_col88[18] <= fa_s0_c88_n601_s;
                    stage1_col88[19] <= fa_s0_c88_n602_s;
                    stage1_col88[20] <= fa_s0_c88_n603_s;
                    stage1_col89[0] <= fa_s0_c88_n593_c;
                    stage1_col89[1] <= fa_s0_c88_n594_c;
                    stage1_col89[2] <= fa_s0_c88_n595_c;
                    stage1_col89[3] <= fa_s0_c88_n596_c;
                    stage1_col89[4] <= fa_s0_c88_n597_c;
                    stage1_col89[5] <= fa_s0_c88_n598_c;
                    stage1_col89[6] <= fa_s0_c88_n599_c;
                    stage1_col89[7] <= fa_s0_c88_n600_c;
                    stage1_col89[8] <= fa_s0_c88_n601_c;
                    stage1_col89[9] <= fa_s0_c88_n602_c;
                    stage1_col89[10] <= fa_s0_c88_n603_c;
                    stage1_col89[11] <= fa_s0_c89_n604_s;
                    stage1_col89[12] <= fa_s0_c89_n605_s;
                    stage1_col89[13] <= fa_s0_c89_n606_s;
                    stage1_col89[14] <= fa_s0_c89_n607_s;
                    stage1_col89[15] <= fa_s0_c89_n608_s;
                    stage1_col89[16] <= fa_s0_c89_n609_s;
                    stage1_col89[17] <= fa_s0_c89_n610_s;
                    stage1_col89[18] <= fa_s0_c89_n611_s;
                    stage1_col89[19] <= fa_s0_c89_n612_s;
                    stage1_col89[20] <= fa_s0_c89_n613_s;
                    stage1_col89[21] <= stage0_col89[30];
                    stage1_col89[22] <= stage0_col89[31];
                    stage1_col90[0] <= fa_s0_c89_n604_c;
                    stage1_col90[1] <= fa_s0_c89_n605_c;
                    stage1_col90[2] <= fa_s0_c89_n606_c;
                    stage1_col90[3] <= fa_s0_c89_n607_c;
                    stage1_col90[4] <= fa_s0_c89_n608_c;
                    stage1_col90[5] <= fa_s0_c89_n609_c;
                    stage1_col90[6] <= fa_s0_c89_n610_c;
                    stage1_col90[7] <= fa_s0_c89_n611_c;
                    stage1_col90[8] <= fa_s0_c89_n612_c;
                    stage1_col90[9] <= fa_s0_c89_n613_c;
                    stage1_col90[10] <= fa_s0_c90_n614_s;
                    stage1_col90[11] <= fa_s0_c90_n615_s;
                    stage1_col90[12] <= fa_s0_c90_n616_s;
                    stage1_col90[13] <= fa_s0_c90_n617_s;
                    stage1_col90[14] <= fa_s0_c90_n618_s;
                    stage1_col90[15] <= fa_s0_c90_n619_s;
                    stage1_col90[16] <= fa_s0_c90_n620_s;
                    stage1_col90[17] <= fa_s0_c90_n621_s;
                    stage1_col90[18] <= fa_s0_c90_n622_s;
                    stage1_col90[19] <= fa_s0_c90_n623_s;
                    stage1_col90[20] <= fa_s0_c90_n624_s;
                    stage1_col91[0] <= fa_s0_c90_n614_c;
                    stage1_col91[1] <= fa_s0_c90_n615_c;
                    stage1_col91[2] <= fa_s0_c90_n616_c;
                    stage1_col91[3] <= fa_s0_c90_n617_c;
                    stage1_col91[4] <= fa_s0_c90_n618_c;
                    stage1_col91[5] <= fa_s0_c90_n619_c;
                    stage1_col91[6] <= fa_s0_c90_n620_c;
                    stage1_col91[7] <= fa_s0_c90_n621_c;
                    stage1_col91[8] <= fa_s0_c90_n622_c;
                    stage1_col91[9] <= fa_s0_c90_n623_c;
                    stage1_col91[10] <= fa_s0_c90_n624_c;
                    stage1_col91[11] <= fa_s0_c91_n625_s;
                    stage1_col91[12] <= fa_s0_c91_n626_s;
                    stage1_col91[13] <= fa_s0_c91_n627_s;
                    stage1_col91[14] <= fa_s0_c91_n628_s;
                    stage1_col91[15] <= fa_s0_c91_n629_s;
                    stage1_col91[16] <= fa_s0_c91_n630_s;
                    stage1_col91[17] <= fa_s0_c91_n631_s;
                    stage1_col91[18] <= fa_s0_c91_n632_s;
                    stage1_col91[19] <= fa_s0_c91_n633_s;
                    stage1_col91[20] <= fa_s0_c91_n634_s;
                    stage1_col91[21] <= stage0_col91[30];
                    stage1_col91[22] <= stage0_col91[31];
                    stage1_col92[0] <= fa_s0_c91_n625_c;
                    stage1_col92[1] <= fa_s0_c91_n626_c;
                    stage1_col92[2] <= fa_s0_c91_n627_c;
                    stage1_col92[3] <= fa_s0_c91_n628_c;
                    stage1_col92[4] <= fa_s0_c91_n629_c;
                    stage1_col92[5] <= fa_s0_c91_n630_c;
                    stage1_col92[6] <= fa_s0_c91_n631_c;
                    stage1_col92[7] <= fa_s0_c91_n632_c;
                    stage1_col92[8] <= fa_s0_c91_n633_c;
                    stage1_col92[9] <= fa_s0_c91_n634_c;
                    stage1_col92[10] <= fa_s0_c92_n635_s;
                    stage1_col92[11] <= fa_s0_c92_n636_s;
                    stage1_col92[12] <= fa_s0_c92_n637_s;
                    stage1_col92[13] <= fa_s0_c92_n638_s;
                    stage1_col92[14] <= fa_s0_c92_n639_s;
                    stage1_col92[15] <= fa_s0_c92_n640_s;
                    stage1_col92[16] <= fa_s0_c92_n641_s;
                    stage1_col92[17] <= fa_s0_c92_n642_s;
                    stage1_col92[18] <= fa_s0_c92_n643_s;
                    stage1_col92[19] <= fa_s0_c92_n644_s;
                    stage1_col92[20] <= fa_s0_c92_n645_s;
                    stage1_col93[0] <= fa_s0_c92_n635_c;
                    stage1_col93[1] <= fa_s0_c92_n636_c;
                    stage1_col93[2] <= fa_s0_c92_n637_c;
                    stage1_col93[3] <= fa_s0_c92_n638_c;
                    stage1_col93[4] <= fa_s0_c92_n639_c;
                    stage1_col93[5] <= fa_s0_c92_n640_c;
                    stage1_col93[6] <= fa_s0_c92_n641_c;
                    stage1_col93[7] <= fa_s0_c92_n642_c;
                    stage1_col93[8] <= fa_s0_c92_n643_c;
                    stage1_col93[9] <= fa_s0_c92_n644_c;
                    stage1_col93[10] <= fa_s0_c92_n645_c;
                    stage1_col93[11] <= fa_s0_c93_n646_s;
                    stage1_col93[12] <= fa_s0_c93_n647_s;
                    stage1_col93[13] <= fa_s0_c93_n648_s;
                    stage1_col93[14] <= fa_s0_c93_n649_s;
                    stage1_col93[15] <= fa_s0_c93_n650_s;
                    stage1_col93[16] <= fa_s0_c93_n651_s;
                    stage1_col93[17] <= fa_s0_c93_n652_s;
                    stage1_col93[18] <= fa_s0_c93_n653_s;
                    stage1_col93[19] <= fa_s0_c93_n654_s;
                    stage1_col93[20] <= fa_s0_c93_n655_s;
                    stage1_col93[21] <= stage0_col93[30];
                    stage1_col93[22] <= stage0_col93[31];
                    stage1_col94[0] <= fa_s0_c93_n646_c;
                    stage1_col94[1] <= fa_s0_c93_n647_c;
                    stage1_col94[2] <= fa_s0_c93_n648_c;
                    stage1_col94[3] <= fa_s0_c93_n649_c;
                    stage1_col94[4] <= fa_s0_c93_n650_c;
                    stage1_col94[5] <= fa_s0_c93_n651_c;
                    stage1_col94[6] <= fa_s0_c93_n652_c;
                    stage1_col94[7] <= fa_s0_c93_n653_c;
                    stage1_col94[8] <= fa_s0_c93_n654_c;
                    stage1_col94[9] <= fa_s0_c93_n655_c;
                    stage1_col94[10] <= fa_s0_c94_n656_s;
                    stage1_col94[11] <= fa_s0_c94_n657_s;
                    stage1_col94[12] <= fa_s0_c94_n658_s;
                    stage1_col94[13] <= fa_s0_c94_n659_s;
                    stage1_col94[14] <= fa_s0_c94_n660_s;
                    stage1_col94[15] <= fa_s0_c94_n661_s;
                    stage1_col94[16] <= fa_s0_c94_n662_s;
                    stage1_col94[17] <= fa_s0_c94_n663_s;
                    stage1_col94[18] <= fa_s0_c94_n664_s;
                    stage1_col94[19] <= fa_s0_c94_n665_s;
                    stage1_col94[20] <= fa_s0_c94_n666_s;
                    stage1_col95[0] <= fa_s0_c94_n656_c;
                    stage1_col95[1] <= fa_s0_c94_n657_c;
                    stage1_col95[2] <= fa_s0_c94_n658_c;
                    stage1_col95[3] <= fa_s0_c94_n659_c;
                    stage1_col95[4] <= fa_s0_c94_n660_c;
                    stage1_col95[5] <= fa_s0_c94_n661_c;
                    stage1_col95[6] <= fa_s0_c94_n662_c;
                    stage1_col95[7] <= fa_s0_c94_n663_c;
                    stage1_col95[8] <= fa_s0_c94_n664_c;
                    stage1_col95[9] <= fa_s0_c94_n665_c;
                    stage1_col95[10] <= fa_s0_c94_n666_c;
                    stage1_col95[11] <= fa_s0_c95_n667_s;
                    stage1_col95[12] <= fa_s0_c95_n668_s;
                    stage1_col95[13] <= fa_s0_c95_n669_s;
                    stage1_col95[14] <= fa_s0_c95_n670_s;
                    stage1_col95[15] <= fa_s0_c95_n671_s;
                    stage1_col95[16] <= fa_s0_c95_n672_s;
                    stage1_col95[17] <= fa_s0_c95_n673_s;
                    stage1_col95[18] <= fa_s0_c95_n674_s;
                    stage1_col95[19] <= fa_s0_c95_n675_s;
                    stage1_col95[20] <= fa_s0_c95_n676_s;
                    stage1_col95[21] <= stage0_col95[30];
                    stage1_col95[22] <= stage0_col95[31];
                    stage1_col96[0] <= fa_s0_c95_n667_c;
                    stage1_col96[1] <= fa_s0_c95_n668_c;
                    stage1_col96[2] <= fa_s0_c95_n669_c;
                    stage1_col96[3] <= fa_s0_c95_n670_c;
                    stage1_col96[4] <= fa_s0_c95_n671_c;
                    stage1_col96[5] <= fa_s0_c95_n672_c;
                    stage1_col96[6] <= fa_s0_c95_n673_c;
                    stage1_col96[7] <= fa_s0_c95_n674_c;
                    stage1_col96[8] <= fa_s0_c95_n675_c;
                    stage1_col96[9] <= fa_s0_c95_n676_c;
                    stage1_col96[10] <= fa_s0_c96_n677_s;
                    stage1_col96[11] <= fa_s0_c96_n678_s;
                    stage1_col96[12] <= fa_s0_c96_n679_s;
                    stage1_col96[13] <= fa_s0_c96_n680_s;
                    stage1_col96[14] <= fa_s0_c96_n681_s;
                    stage1_col96[15] <= fa_s0_c96_n682_s;
                    stage1_col96[16] <= fa_s0_c96_n683_s;
                    stage1_col96[17] <= fa_s0_c96_n684_s;
                    stage1_col96[18] <= fa_s0_c96_n685_s;
                    stage1_col96[19] <= fa_s0_c96_n686_s;
                    stage1_col96[20] <= fa_s0_c96_n687_s;
                    stage1_col97[0] <= fa_s0_c96_n677_c;
                    stage1_col97[1] <= fa_s0_c96_n678_c;
                    stage1_col97[2] <= fa_s0_c96_n679_c;
                    stage1_col97[3] <= fa_s0_c96_n680_c;
                    stage1_col97[4] <= fa_s0_c96_n681_c;
                    stage1_col97[5] <= fa_s0_c96_n682_c;
                    stage1_col97[6] <= fa_s0_c96_n683_c;
                    stage1_col97[7] <= fa_s0_c96_n684_c;
                    stage1_col97[8] <= fa_s0_c96_n685_c;
                    stage1_col97[9] <= fa_s0_c96_n686_c;
                    stage1_col97[10] <= fa_s0_c96_n687_c;
                    stage1_col97[11] <= fa_s0_c97_n688_s;
                    stage1_col97[12] <= fa_s0_c97_n689_s;
                    stage1_col97[13] <= fa_s0_c97_n690_s;
                    stage1_col97[14] <= fa_s0_c97_n691_s;
                    stage1_col97[15] <= fa_s0_c97_n692_s;
                    stage1_col97[16] <= fa_s0_c97_n693_s;
                    stage1_col97[17] <= fa_s0_c97_n694_s;
                    stage1_col97[18] <= fa_s0_c97_n695_s;
                    stage1_col97[19] <= fa_s0_c97_n696_s;
                    stage1_col97[20] <= fa_s0_c97_n697_s;
                    stage1_col97[21] <= stage0_col97[30];
                    stage1_col97[22] <= stage0_col97[31];
                    stage1_col98[0] <= fa_s0_c97_n688_c;
                    stage1_col98[1] <= fa_s0_c97_n689_c;
                    stage1_col98[2] <= fa_s0_c97_n690_c;
                    stage1_col98[3] <= fa_s0_c97_n691_c;
                    stage1_col98[4] <= fa_s0_c97_n692_c;
                    stage1_col98[5] <= fa_s0_c97_n693_c;
                    stage1_col98[6] <= fa_s0_c97_n694_c;
                    stage1_col98[7] <= fa_s0_c97_n695_c;
                    stage1_col98[8] <= fa_s0_c97_n696_c;
                    stage1_col98[9] <= fa_s0_c97_n697_c;
                    stage1_col98[10] <= fa_s0_c98_n698_s;
                    stage1_col98[11] <= fa_s0_c98_n699_s;
                    stage1_col98[12] <= fa_s0_c98_n700_s;
                    stage1_col98[13] <= fa_s0_c98_n701_s;
                    stage1_col98[14] <= fa_s0_c98_n702_s;
                    stage1_col98[15] <= fa_s0_c98_n703_s;
                    stage1_col98[16] <= fa_s0_c98_n704_s;
                    stage1_col98[17] <= fa_s0_c98_n705_s;
                    stage1_col98[18] <= fa_s0_c98_n706_s;
                    stage1_col98[19] <= fa_s0_c98_n707_s;
                    stage1_col98[20] <= fa_s0_c98_n708_s;
                    stage1_col99[0] <= fa_s0_c98_n698_c;
                    stage1_col99[1] <= fa_s0_c98_n699_c;
                    stage1_col99[2] <= fa_s0_c98_n700_c;
                    stage1_col99[3] <= fa_s0_c98_n701_c;
                    stage1_col99[4] <= fa_s0_c98_n702_c;
                    stage1_col99[5] <= fa_s0_c98_n703_c;
                    stage1_col99[6] <= fa_s0_c98_n704_c;
                    stage1_col99[7] <= fa_s0_c98_n705_c;
                    stage1_col99[8] <= fa_s0_c98_n706_c;
                    stage1_col99[9] <= fa_s0_c98_n707_c;
                    stage1_col99[10] <= fa_s0_c98_n708_c;
                    stage1_col99[11] <= fa_s0_c99_n709_s;
                    stage1_col99[12] <= fa_s0_c99_n710_s;
                    stage1_col99[13] <= fa_s0_c99_n711_s;
                    stage1_col99[14] <= fa_s0_c99_n712_s;
                    stage1_col99[15] <= fa_s0_c99_n713_s;
                    stage1_col99[16] <= fa_s0_c99_n714_s;
                    stage1_col99[17] <= fa_s0_c99_n715_s;
                    stage1_col99[18] <= fa_s0_c99_n716_s;
                    stage1_col99[19] <= fa_s0_c99_n717_s;
                    stage1_col99[20] <= fa_s0_c99_n718_s;
                    stage1_col99[21] <= stage0_col99[30];
                    stage1_col99[22] <= stage0_col99[31];
                    stage1_col100[0] <= fa_s0_c99_n709_c;
                    stage1_col100[1] <= fa_s0_c99_n710_c;
                    stage1_col100[2] <= fa_s0_c99_n711_c;
                    stage1_col100[3] <= fa_s0_c99_n712_c;
                    stage1_col100[4] <= fa_s0_c99_n713_c;
                    stage1_col100[5] <= fa_s0_c99_n714_c;
                    stage1_col100[6] <= fa_s0_c99_n715_c;
                    stage1_col100[7] <= fa_s0_c99_n716_c;
                    stage1_col100[8] <= fa_s0_c99_n717_c;
                    stage1_col100[9] <= fa_s0_c99_n718_c;
                    stage1_col100[10] <= fa_s0_c100_n719_s;
                    stage1_col100[11] <= fa_s0_c100_n720_s;
                    stage1_col100[12] <= fa_s0_c100_n721_s;
                    stage1_col100[13] <= fa_s0_c100_n722_s;
                    stage1_col100[14] <= fa_s0_c100_n723_s;
                    stage1_col100[15] <= fa_s0_c100_n724_s;
                    stage1_col100[16] <= fa_s0_c100_n725_s;
                    stage1_col100[17] <= fa_s0_c100_n726_s;
                    stage1_col100[18] <= fa_s0_c100_n727_s;
                    stage1_col100[19] <= fa_s0_c100_n728_s;
                    stage1_col100[20] <= fa_s0_c100_n729_s;
                    stage1_col101[0] <= fa_s0_c100_n719_c;
                    stage1_col101[1] <= fa_s0_c100_n720_c;
                    stage1_col101[2] <= fa_s0_c100_n721_c;
                    stage1_col101[3] <= fa_s0_c100_n722_c;
                    stage1_col101[4] <= fa_s0_c100_n723_c;
                    stage1_col101[5] <= fa_s0_c100_n724_c;
                    stage1_col101[6] <= fa_s0_c100_n725_c;
                    stage1_col101[7] <= fa_s0_c100_n726_c;
                    stage1_col101[8] <= fa_s0_c100_n727_c;
                    stage1_col101[9] <= fa_s0_c100_n728_c;
                    stage1_col101[10] <= fa_s0_c100_n729_c;
                    stage1_col101[11] <= fa_s0_c101_n730_s;
                    stage1_col101[12] <= fa_s0_c101_n731_s;
                    stage1_col101[13] <= fa_s0_c101_n732_s;
                    stage1_col101[14] <= fa_s0_c101_n733_s;
                    stage1_col101[15] <= fa_s0_c101_n734_s;
                    stage1_col101[16] <= fa_s0_c101_n735_s;
                    stage1_col101[17] <= fa_s0_c101_n736_s;
                    stage1_col101[18] <= fa_s0_c101_n737_s;
                    stage1_col101[19] <= fa_s0_c101_n738_s;
                    stage1_col101[20] <= fa_s0_c101_n739_s;
                    stage1_col101[21] <= stage0_col101[30];
                    stage1_col101[22] <= stage0_col101[31];
                    stage1_col102[0] <= fa_s0_c101_n730_c;
                    stage1_col102[1] <= fa_s0_c101_n731_c;
                    stage1_col102[2] <= fa_s0_c101_n732_c;
                    stage1_col102[3] <= fa_s0_c101_n733_c;
                    stage1_col102[4] <= fa_s0_c101_n734_c;
                    stage1_col102[5] <= fa_s0_c101_n735_c;
                    stage1_col102[6] <= fa_s0_c101_n736_c;
                    stage1_col102[7] <= fa_s0_c101_n737_c;
                    stage1_col102[8] <= fa_s0_c101_n738_c;
                    stage1_col102[9] <= fa_s0_c101_n739_c;
                    stage1_col102[10] <= fa_s0_c102_n740_s;
                    stage1_col102[11] <= fa_s0_c102_n741_s;
                    stage1_col102[12] <= fa_s0_c102_n742_s;
                    stage1_col102[13] <= fa_s0_c102_n743_s;
                    stage1_col102[14] <= fa_s0_c102_n744_s;
                    stage1_col102[15] <= fa_s0_c102_n745_s;
                    stage1_col102[16] <= fa_s0_c102_n746_s;
                    stage1_col102[17] <= fa_s0_c102_n747_s;
                    stage1_col102[18] <= fa_s0_c102_n748_s;
                    stage1_col102[19] <= fa_s0_c102_n749_s;
                    stage1_col102[20] <= fa_s0_c102_n750_s;
                    stage1_col103[0] <= fa_s0_c102_n740_c;
                    stage1_col103[1] <= fa_s0_c102_n741_c;
                    stage1_col103[2] <= fa_s0_c102_n742_c;
                    stage1_col103[3] <= fa_s0_c102_n743_c;
                    stage1_col103[4] <= fa_s0_c102_n744_c;
                    stage1_col103[5] <= fa_s0_c102_n745_c;
                    stage1_col103[6] <= fa_s0_c102_n746_c;
                    stage1_col103[7] <= fa_s0_c102_n747_c;
                    stage1_col103[8] <= fa_s0_c102_n748_c;
                    stage1_col103[9] <= fa_s0_c102_n749_c;
                    stage1_col103[10] <= fa_s0_c102_n750_c;
                    stage1_col103[11] <= fa_s0_c103_n751_s;
                    stage1_col103[12] <= fa_s0_c103_n752_s;
                    stage1_col103[13] <= fa_s0_c103_n753_s;
                    stage1_col103[14] <= fa_s0_c103_n754_s;
                    stage1_col103[15] <= fa_s0_c103_n755_s;
                    stage1_col103[16] <= fa_s0_c103_n756_s;
                    stage1_col103[17] <= fa_s0_c103_n757_s;
                    stage1_col103[18] <= fa_s0_c103_n758_s;
                    stage1_col103[19] <= fa_s0_c103_n759_s;
                    stage1_col103[20] <= fa_s0_c103_n760_s;
                    stage1_col103[21] <= stage0_col103[30];
                    stage1_col103[22] <= stage0_col103[31];
                    stage1_col104[0] <= fa_s0_c103_n751_c;
                    stage1_col104[1] <= fa_s0_c103_n752_c;
                    stage1_col104[2] <= fa_s0_c103_n753_c;
                    stage1_col104[3] <= fa_s0_c103_n754_c;
                    stage1_col104[4] <= fa_s0_c103_n755_c;
                    stage1_col104[5] <= fa_s0_c103_n756_c;
                    stage1_col104[6] <= fa_s0_c103_n757_c;
                    stage1_col104[7] <= fa_s0_c103_n758_c;
                    stage1_col104[8] <= fa_s0_c103_n759_c;
                    stage1_col104[9] <= fa_s0_c103_n760_c;
                    stage1_col104[10] <= fa_s0_c104_n761_s;
                    stage1_col104[11] <= fa_s0_c104_n762_s;
                    stage1_col104[12] <= fa_s0_c104_n763_s;
                    stage1_col104[13] <= fa_s0_c104_n764_s;
                    stage1_col104[14] <= fa_s0_c104_n765_s;
                    stage1_col104[15] <= fa_s0_c104_n766_s;
                    stage1_col104[16] <= fa_s0_c104_n767_s;
                    stage1_col104[17] <= fa_s0_c104_n768_s;
                    stage1_col104[18] <= fa_s0_c104_n769_s;
                    stage1_col104[19] <= fa_s0_c104_n770_s;
                    stage1_col104[20] <= fa_s0_c104_n771_s;
                    stage1_col105[0] <= fa_s0_c104_n761_c;
                    stage1_col105[1] <= fa_s0_c104_n762_c;
                    stage1_col105[2] <= fa_s0_c104_n763_c;
                    stage1_col105[3] <= fa_s0_c104_n764_c;
                    stage1_col105[4] <= fa_s0_c104_n765_c;
                    stage1_col105[5] <= fa_s0_c104_n766_c;
                    stage1_col105[6] <= fa_s0_c104_n767_c;
                    stage1_col105[7] <= fa_s0_c104_n768_c;
                    stage1_col105[8] <= fa_s0_c104_n769_c;
                    stage1_col105[9] <= fa_s0_c104_n770_c;
                    stage1_col105[10] <= fa_s0_c104_n771_c;
                    stage1_col105[11] <= fa_s0_c105_n772_s;
                    stage1_col105[12] <= fa_s0_c105_n773_s;
                    stage1_col105[13] <= fa_s0_c105_n774_s;
                    stage1_col105[14] <= fa_s0_c105_n775_s;
                    stage1_col105[15] <= fa_s0_c105_n776_s;
                    stage1_col105[16] <= fa_s0_c105_n777_s;
                    stage1_col105[17] <= fa_s0_c105_n778_s;
                    stage1_col105[18] <= fa_s0_c105_n779_s;
                    stage1_col105[19] <= fa_s0_c105_n780_s;
                    stage1_col105[20] <= fa_s0_c105_n781_s;
                    stage1_col105[21] <= stage0_col105[30];
                    stage1_col105[22] <= stage0_col105[31];
                    stage1_col106[0] <= fa_s0_c105_n772_c;
                    stage1_col106[1] <= fa_s0_c105_n773_c;
                    stage1_col106[2] <= fa_s0_c105_n774_c;
                    stage1_col106[3] <= fa_s0_c105_n775_c;
                    stage1_col106[4] <= fa_s0_c105_n776_c;
                    stage1_col106[5] <= fa_s0_c105_n777_c;
                    stage1_col106[6] <= fa_s0_c105_n778_c;
                    stage1_col106[7] <= fa_s0_c105_n779_c;
                    stage1_col106[8] <= fa_s0_c105_n780_c;
                    stage1_col106[9] <= fa_s0_c105_n781_c;
                    stage1_col106[10] <= fa_s0_c106_n782_s;
                    stage1_col106[11] <= fa_s0_c106_n783_s;
                    stage1_col106[12] <= fa_s0_c106_n784_s;
                    stage1_col106[13] <= fa_s0_c106_n785_s;
                    stage1_col106[14] <= fa_s0_c106_n786_s;
                    stage1_col106[15] <= fa_s0_c106_n787_s;
                    stage1_col106[16] <= fa_s0_c106_n788_s;
                    stage1_col106[17] <= fa_s0_c106_n789_s;
                    stage1_col106[18] <= fa_s0_c106_n790_s;
                    stage1_col106[19] <= fa_s0_c106_n791_s;
                    stage1_col106[20] <= fa_s0_c106_n792_s;
                    stage1_col107[0] <= fa_s0_c106_n782_c;
                    stage1_col107[1] <= fa_s0_c106_n783_c;
                    stage1_col107[2] <= fa_s0_c106_n784_c;
                    stage1_col107[3] <= fa_s0_c106_n785_c;
                    stage1_col107[4] <= fa_s0_c106_n786_c;
                    stage1_col107[5] <= fa_s0_c106_n787_c;
                    stage1_col107[6] <= fa_s0_c106_n788_c;
                    stage1_col107[7] <= fa_s0_c106_n789_c;
                    stage1_col107[8] <= fa_s0_c106_n790_c;
                    stage1_col107[9] <= fa_s0_c106_n791_c;
                    stage1_col107[10] <= fa_s0_c106_n792_c;
                    stage1_col107[11] <= fa_s0_c107_n793_s;
                    stage1_col107[12] <= fa_s0_c107_n794_s;
                    stage1_col107[13] <= fa_s0_c107_n795_s;
                    stage1_col107[14] <= fa_s0_c107_n796_s;
                    stage1_col107[15] <= fa_s0_c107_n797_s;
                    stage1_col107[16] <= fa_s0_c107_n798_s;
                    stage1_col107[17] <= fa_s0_c107_n799_s;
                    stage1_col107[18] <= fa_s0_c107_n800_s;
                    stage1_col107[19] <= fa_s0_c107_n801_s;
                    stage1_col107[20] <= fa_s0_c107_n802_s;
                    stage1_col107[21] <= stage0_col107[30];
                    stage1_col107[22] <= stage0_col107[31];
                    stage1_col108[0] <= fa_s0_c107_n793_c;
                    stage1_col108[1] <= fa_s0_c107_n794_c;
                    stage1_col108[2] <= fa_s0_c107_n795_c;
                    stage1_col108[3] <= fa_s0_c107_n796_c;
                    stage1_col108[4] <= fa_s0_c107_n797_c;
                    stage1_col108[5] <= fa_s0_c107_n798_c;
                    stage1_col108[6] <= fa_s0_c107_n799_c;
                    stage1_col108[7] <= fa_s0_c107_n800_c;
                    stage1_col108[8] <= fa_s0_c107_n801_c;
                    stage1_col108[9] <= fa_s0_c107_n802_c;
                    stage1_col108[10] <= fa_s0_c108_n803_s;
                    stage1_col108[11] <= fa_s0_c108_n804_s;
                    stage1_col108[12] <= fa_s0_c108_n805_s;
                    stage1_col108[13] <= fa_s0_c108_n806_s;
                    stage1_col108[14] <= fa_s0_c108_n807_s;
                    stage1_col108[15] <= fa_s0_c108_n808_s;
                    stage1_col108[16] <= fa_s0_c108_n809_s;
                    stage1_col108[17] <= fa_s0_c108_n810_s;
                    stage1_col108[18] <= fa_s0_c108_n811_s;
                    stage1_col108[19] <= fa_s0_c108_n812_s;
                    stage1_col108[20] <= fa_s0_c108_n813_s;
                    stage1_col109[0] <= fa_s0_c108_n803_c;
                    stage1_col109[1] <= fa_s0_c108_n804_c;
                    stage1_col109[2] <= fa_s0_c108_n805_c;
                    stage1_col109[3] <= fa_s0_c108_n806_c;
                    stage1_col109[4] <= fa_s0_c108_n807_c;
                    stage1_col109[5] <= fa_s0_c108_n808_c;
                    stage1_col109[6] <= fa_s0_c108_n809_c;
                    stage1_col109[7] <= fa_s0_c108_n810_c;
                    stage1_col109[8] <= fa_s0_c108_n811_c;
                    stage1_col109[9] <= fa_s0_c108_n812_c;
                    stage1_col109[10] <= fa_s0_c108_n813_c;
                    stage1_col109[11] <= fa_s0_c109_n814_s;
                    stage1_col109[12] <= fa_s0_c109_n815_s;
                    stage1_col109[13] <= fa_s0_c109_n816_s;
                    stage1_col109[14] <= fa_s0_c109_n817_s;
                    stage1_col109[15] <= fa_s0_c109_n818_s;
                    stage1_col109[16] <= fa_s0_c109_n819_s;
                    stage1_col109[17] <= fa_s0_c109_n820_s;
                    stage1_col109[18] <= fa_s0_c109_n821_s;
                    stage1_col109[19] <= fa_s0_c109_n822_s;
                    stage1_col109[20] <= fa_s0_c109_n823_s;
                    stage1_col109[21] <= stage0_col109[30];
                    stage1_col109[22] <= stage0_col109[31];
                    stage1_col110[0] <= fa_s0_c109_n814_c;
                    stage1_col110[1] <= fa_s0_c109_n815_c;
                    stage1_col110[2] <= fa_s0_c109_n816_c;
                    stage1_col110[3] <= fa_s0_c109_n817_c;
                    stage1_col110[4] <= fa_s0_c109_n818_c;
                    stage1_col110[5] <= fa_s0_c109_n819_c;
                    stage1_col110[6] <= fa_s0_c109_n820_c;
                    stage1_col110[7] <= fa_s0_c109_n821_c;
                    stage1_col110[8] <= fa_s0_c109_n822_c;
                    stage1_col110[9] <= fa_s0_c109_n823_c;
                    stage1_col110[10] <= fa_s0_c110_n824_s;
                    stage1_col110[11] <= fa_s0_c110_n825_s;
                    stage1_col110[12] <= fa_s0_c110_n826_s;
                    stage1_col110[13] <= fa_s0_c110_n827_s;
                    stage1_col110[14] <= fa_s0_c110_n828_s;
                    stage1_col110[15] <= fa_s0_c110_n829_s;
                    stage1_col110[16] <= fa_s0_c110_n830_s;
                    stage1_col110[17] <= fa_s0_c110_n831_s;
                    stage1_col110[18] <= fa_s0_c110_n832_s;
                    stage1_col110[19] <= fa_s0_c110_n833_s;
                    stage1_col110[20] <= fa_s0_c110_n834_s;
                    stage1_col111[0] <= fa_s0_c110_n824_c;
                    stage1_col111[1] <= fa_s0_c110_n825_c;
                    stage1_col111[2] <= fa_s0_c110_n826_c;
                    stage1_col111[3] <= fa_s0_c110_n827_c;
                    stage1_col111[4] <= fa_s0_c110_n828_c;
                    stage1_col111[5] <= fa_s0_c110_n829_c;
                    stage1_col111[6] <= fa_s0_c110_n830_c;
                    stage1_col111[7] <= fa_s0_c110_n831_c;
                    stage1_col111[8] <= fa_s0_c110_n832_c;
                    stage1_col111[9] <= fa_s0_c110_n833_c;
                    stage1_col111[10] <= fa_s0_c110_n834_c;
                    stage1_col111[11] <= fa_s0_c111_n835_s;
                    stage1_col111[12] <= fa_s0_c111_n836_s;
                    stage1_col111[13] <= fa_s0_c111_n837_s;
                    stage1_col111[14] <= fa_s0_c111_n838_s;
                    stage1_col111[15] <= fa_s0_c111_n839_s;
                    stage1_col111[16] <= fa_s0_c111_n840_s;
                    stage1_col111[17] <= fa_s0_c111_n841_s;
                    stage1_col111[18] <= fa_s0_c111_n842_s;
                    stage1_col111[19] <= fa_s0_c111_n843_s;
                    stage1_col111[20] <= fa_s0_c111_n844_s;
                    stage1_col111[21] <= stage0_col111[30];
                    stage1_col111[22] <= stage0_col111[31];
                    stage1_col112[0] <= fa_s0_c111_n835_c;
                    stage1_col112[1] <= fa_s0_c111_n836_c;
                    stage1_col112[2] <= fa_s0_c111_n837_c;
                    stage1_col112[3] <= fa_s0_c111_n838_c;
                    stage1_col112[4] <= fa_s0_c111_n839_c;
                    stage1_col112[5] <= fa_s0_c111_n840_c;
                    stage1_col112[6] <= fa_s0_c111_n841_c;
                    stage1_col112[7] <= fa_s0_c111_n842_c;
                    stage1_col112[8] <= fa_s0_c111_n843_c;
                    stage1_col112[9] <= fa_s0_c111_n844_c;
                    stage1_col112[10] <= fa_s0_c112_n845_s;
                    stage1_col112[11] <= fa_s0_c112_n846_s;
                    stage1_col112[12] <= fa_s0_c112_n847_s;
                    stage1_col112[13] <= fa_s0_c112_n848_s;
                    stage1_col112[14] <= fa_s0_c112_n849_s;
                    stage1_col112[15] <= fa_s0_c112_n850_s;
                    stage1_col112[16] <= fa_s0_c112_n851_s;
                    stage1_col112[17] <= fa_s0_c112_n852_s;
                    stage1_col112[18] <= fa_s0_c112_n853_s;
                    stage1_col112[19] <= fa_s0_c112_n854_s;
                    stage1_col112[20] <= fa_s0_c112_n855_s;
                    stage1_col113[0] <= fa_s0_c112_n845_c;
                    stage1_col113[1] <= fa_s0_c112_n846_c;
                    stage1_col113[2] <= fa_s0_c112_n847_c;
                    stage1_col113[3] <= fa_s0_c112_n848_c;
                    stage1_col113[4] <= fa_s0_c112_n849_c;
                    stage1_col113[5] <= fa_s0_c112_n850_c;
                    stage1_col113[6] <= fa_s0_c112_n851_c;
                    stage1_col113[7] <= fa_s0_c112_n852_c;
                    stage1_col113[8] <= fa_s0_c112_n853_c;
                    stage1_col113[9] <= fa_s0_c112_n854_c;
                    stage1_col113[10] <= fa_s0_c112_n855_c;
                    stage1_col113[11] <= fa_s0_c113_n856_s;
                    stage1_col113[12] <= fa_s0_c113_n857_s;
                    stage1_col113[13] <= fa_s0_c113_n858_s;
                    stage1_col113[14] <= fa_s0_c113_n859_s;
                    stage1_col113[15] <= fa_s0_c113_n860_s;
                    stage1_col113[16] <= fa_s0_c113_n861_s;
                    stage1_col113[17] <= fa_s0_c113_n862_s;
                    stage1_col113[18] <= fa_s0_c113_n863_s;
                    stage1_col113[19] <= fa_s0_c113_n864_s;
                    stage1_col113[20] <= fa_s0_c113_n865_s;
                    stage1_col113[21] <= stage0_col113[30];
                    stage1_col113[22] <= stage0_col113[31];
                    stage1_col114[0] <= fa_s0_c113_n856_c;
                    stage1_col114[1] <= fa_s0_c113_n857_c;
                    stage1_col114[2] <= fa_s0_c113_n858_c;
                    stage1_col114[3] <= fa_s0_c113_n859_c;
                    stage1_col114[4] <= fa_s0_c113_n860_c;
                    stage1_col114[5] <= fa_s0_c113_n861_c;
                    stage1_col114[6] <= fa_s0_c113_n862_c;
                    stage1_col114[7] <= fa_s0_c113_n863_c;
                    stage1_col114[8] <= fa_s0_c113_n864_c;
                    stage1_col114[9] <= fa_s0_c113_n865_c;
                    stage1_col114[10] <= fa_s0_c114_n866_s;
                    stage1_col114[11] <= fa_s0_c114_n867_s;
                    stage1_col114[12] <= fa_s0_c114_n868_s;
                    stage1_col114[13] <= fa_s0_c114_n869_s;
                    stage1_col114[14] <= fa_s0_c114_n870_s;
                    stage1_col114[15] <= fa_s0_c114_n871_s;
                    stage1_col114[16] <= fa_s0_c114_n872_s;
                    stage1_col114[17] <= fa_s0_c114_n873_s;
                    stage1_col114[18] <= fa_s0_c114_n874_s;
                    stage1_col114[19] <= fa_s0_c114_n875_s;
                    stage1_col114[20] <= fa_s0_c114_n876_s;
                    stage1_col115[0] <= fa_s0_c114_n866_c;
                    stage1_col115[1] <= fa_s0_c114_n867_c;
                    stage1_col115[2] <= fa_s0_c114_n868_c;
                    stage1_col115[3] <= fa_s0_c114_n869_c;
                    stage1_col115[4] <= fa_s0_c114_n870_c;
                    stage1_col115[5] <= fa_s0_c114_n871_c;
                    stage1_col115[6] <= fa_s0_c114_n872_c;
                    stage1_col115[7] <= fa_s0_c114_n873_c;
                    stage1_col115[8] <= fa_s0_c114_n874_c;
                    stage1_col115[9] <= fa_s0_c114_n875_c;
                    stage1_col115[10] <= fa_s0_c114_n876_c;
                    stage1_col115[11] <= fa_s0_c115_n877_s;
                    stage1_col115[12] <= fa_s0_c115_n878_s;
                    stage1_col115[13] <= fa_s0_c115_n879_s;
                    stage1_col115[14] <= fa_s0_c115_n880_s;
                    stage1_col115[15] <= fa_s0_c115_n881_s;
                    stage1_col115[16] <= fa_s0_c115_n882_s;
                    stage1_col115[17] <= fa_s0_c115_n883_s;
                    stage1_col115[18] <= fa_s0_c115_n884_s;
                    stage1_col115[19] <= fa_s0_c115_n885_s;
                    stage1_col115[20] <= fa_s0_c115_n886_s;
                    stage1_col115[21] <= stage0_col115[30];
                    stage1_col115[22] <= stage0_col115[31];
                    stage1_col116[0] <= fa_s0_c115_n877_c;
                    stage1_col116[1] <= fa_s0_c115_n878_c;
                    stage1_col116[2] <= fa_s0_c115_n879_c;
                    stage1_col116[3] <= fa_s0_c115_n880_c;
                    stage1_col116[4] <= fa_s0_c115_n881_c;
                    stage1_col116[5] <= fa_s0_c115_n882_c;
                    stage1_col116[6] <= fa_s0_c115_n883_c;
                    stage1_col116[7] <= fa_s0_c115_n884_c;
                    stage1_col116[8] <= fa_s0_c115_n885_c;
                    stage1_col116[9] <= fa_s0_c115_n886_c;
                    stage1_col116[10] <= fa_s0_c116_n887_s;
                    stage1_col116[11] <= fa_s0_c116_n888_s;
                    stage1_col116[12] <= fa_s0_c116_n889_s;
                    stage1_col116[13] <= fa_s0_c116_n890_s;
                    stage1_col116[14] <= fa_s0_c116_n891_s;
                    stage1_col116[15] <= fa_s0_c116_n892_s;
                    stage1_col116[16] <= fa_s0_c116_n893_s;
                    stage1_col116[17] <= fa_s0_c116_n894_s;
                    stage1_col116[18] <= fa_s0_c116_n895_s;
                    stage1_col116[19] <= fa_s0_c116_n896_s;
                    stage1_col116[20] <= fa_s0_c116_n897_s;
                    stage1_col117[0] <= fa_s0_c116_n887_c;
                    stage1_col117[1] <= fa_s0_c116_n888_c;
                    stage1_col117[2] <= fa_s0_c116_n889_c;
                    stage1_col117[3] <= fa_s0_c116_n890_c;
                    stage1_col117[4] <= fa_s0_c116_n891_c;
                    stage1_col117[5] <= fa_s0_c116_n892_c;
                    stage1_col117[6] <= fa_s0_c116_n893_c;
                    stage1_col117[7] <= fa_s0_c116_n894_c;
                    stage1_col117[8] <= fa_s0_c116_n895_c;
                    stage1_col117[9] <= fa_s0_c116_n896_c;
                    stage1_col117[10] <= fa_s0_c116_n897_c;
                    stage1_col117[11] <= fa_s0_c117_n898_s;
                    stage1_col117[12] <= fa_s0_c117_n899_s;
                    stage1_col117[13] <= fa_s0_c117_n900_s;
                    stage1_col117[14] <= fa_s0_c117_n901_s;
                    stage1_col117[15] <= fa_s0_c117_n902_s;
                    stage1_col117[16] <= fa_s0_c117_n903_s;
                    stage1_col117[17] <= fa_s0_c117_n904_s;
                    stage1_col117[18] <= fa_s0_c117_n905_s;
                    stage1_col117[19] <= fa_s0_c117_n906_s;
                    stage1_col117[20] <= fa_s0_c117_n907_s;
                    stage1_col117[21] <= stage0_col117[30];
                    stage1_col117[22] <= stage0_col117[31];
                    stage1_col118[0] <= fa_s0_c117_n898_c;
                    stage1_col118[1] <= fa_s0_c117_n899_c;
                    stage1_col118[2] <= fa_s0_c117_n900_c;
                    stage1_col118[3] <= fa_s0_c117_n901_c;
                    stage1_col118[4] <= fa_s0_c117_n902_c;
                    stage1_col118[5] <= fa_s0_c117_n903_c;
                    stage1_col118[6] <= fa_s0_c117_n904_c;
                    stage1_col118[7] <= fa_s0_c117_n905_c;
                    stage1_col118[8] <= fa_s0_c117_n906_c;
                    stage1_col118[9] <= fa_s0_c117_n907_c;
                    stage1_col118[10] <= fa_s0_c118_n908_s;
                    stage1_col118[11] <= fa_s0_c118_n909_s;
                    stage1_col118[12] <= fa_s0_c118_n910_s;
                    stage1_col118[13] <= fa_s0_c118_n911_s;
                    stage1_col118[14] <= fa_s0_c118_n912_s;
                    stage1_col118[15] <= fa_s0_c118_n913_s;
                    stage1_col118[16] <= fa_s0_c118_n914_s;
                    stage1_col118[17] <= fa_s0_c118_n915_s;
                    stage1_col118[18] <= fa_s0_c118_n916_s;
                    stage1_col118[19] <= fa_s0_c118_n917_s;
                    stage1_col118[20] <= fa_s0_c118_n918_s;
                    stage1_col119[0] <= fa_s0_c118_n908_c;
                    stage1_col119[1] <= fa_s0_c118_n909_c;
                    stage1_col119[2] <= fa_s0_c118_n910_c;
                    stage1_col119[3] <= fa_s0_c118_n911_c;
                    stage1_col119[4] <= fa_s0_c118_n912_c;
                    stage1_col119[5] <= fa_s0_c118_n913_c;
                    stage1_col119[6] <= fa_s0_c118_n914_c;
                    stage1_col119[7] <= fa_s0_c118_n915_c;
                    stage1_col119[8] <= fa_s0_c118_n916_c;
                    stage1_col119[9] <= fa_s0_c118_n917_c;
                    stage1_col119[10] <= fa_s0_c118_n918_c;
                    stage1_col119[11] <= fa_s0_c119_n919_s;
                    stage1_col119[12] <= fa_s0_c119_n920_s;
                    stage1_col119[13] <= fa_s0_c119_n921_s;
                    stage1_col119[14] <= fa_s0_c119_n922_s;
                    stage1_col119[15] <= fa_s0_c119_n923_s;
                    stage1_col119[16] <= fa_s0_c119_n924_s;
                    stage1_col119[17] <= fa_s0_c119_n925_s;
                    stage1_col119[18] <= fa_s0_c119_n926_s;
                    stage1_col119[19] <= fa_s0_c119_n927_s;
                    stage1_col119[20] <= fa_s0_c119_n928_s;
                    stage1_col119[21] <= stage0_col119[30];
                    stage1_col119[22] <= stage0_col119[31];
                    stage1_col120[0] <= fa_s0_c119_n919_c;
                    stage1_col120[1] <= fa_s0_c119_n920_c;
                    stage1_col120[2] <= fa_s0_c119_n921_c;
                    stage1_col120[3] <= fa_s0_c119_n922_c;
                    stage1_col120[4] <= fa_s0_c119_n923_c;
                    stage1_col120[5] <= fa_s0_c119_n924_c;
                    stage1_col120[6] <= fa_s0_c119_n925_c;
                    stage1_col120[7] <= fa_s0_c119_n926_c;
                    stage1_col120[8] <= fa_s0_c119_n927_c;
                    stage1_col120[9] <= fa_s0_c119_n928_c;
                    stage1_col120[10] <= fa_s0_c120_n929_s;
                    stage1_col120[11] <= fa_s0_c120_n930_s;
                    stage1_col120[12] <= fa_s0_c120_n931_s;
                    stage1_col120[13] <= fa_s0_c120_n932_s;
                    stage1_col120[14] <= fa_s0_c120_n933_s;
                    stage1_col120[15] <= fa_s0_c120_n934_s;
                    stage1_col120[16] <= fa_s0_c120_n935_s;
                    stage1_col120[17] <= fa_s0_c120_n936_s;
                    stage1_col120[18] <= fa_s0_c120_n937_s;
                    stage1_col120[19] <= fa_s0_c120_n938_s;
                    stage1_col120[20] <= fa_s0_c120_n939_s;
                    stage1_col121[0] <= fa_s0_c120_n929_c;
                    stage1_col121[1] <= fa_s0_c120_n930_c;
                    stage1_col121[2] <= fa_s0_c120_n931_c;
                    stage1_col121[3] <= fa_s0_c120_n932_c;
                    stage1_col121[4] <= fa_s0_c120_n933_c;
                    stage1_col121[5] <= fa_s0_c120_n934_c;
                    stage1_col121[6] <= fa_s0_c120_n935_c;
                    stage1_col121[7] <= fa_s0_c120_n936_c;
                    stage1_col121[8] <= fa_s0_c120_n937_c;
                    stage1_col121[9] <= fa_s0_c120_n938_c;
                    stage1_col121[10] <= fa_s0_c120_n939_c;
                    stage1_col121[11] <= fa_s0_c121_n940_s;
                    stage1_col121[12] <= fa_s0_c121_n941_s;
                    stage1_col121[13] <= fa_s0_c121_n942_s;
                    stage1_col121[14] <= fa_s0_c121_n943_s;
                    stage1_col121[15] <= fa_s0_c121_n944_s;
                    stage1_col121[16] <= fa_s0_c121_n945_s;
                    stage1_col121[17] <= fa_s0_c121_n946_s;
                    stage1_col121[18] <= fa_s0_c121_n947_s;
                    stage1_col121[19] <= fa_s0_c121_n948_s;
                    stage1_col121[20] <= fa_s0_c121_n949_s;
                    stage1_col121[21] <= stage0_col121[30];
                    stage1_col121[22] <= stage0_col121[31];
                    stage1_col122[0] <= fa_s0_c121_n940_c;
                    stage1_col122[1] <= fa_s0_c121_n941_c;
                    stage1_col122[2] <= fa_s0_c121_n942_c;
                    stage1_col122[3] <= fa_s0_c121_n943_c;
                    stage1_col122[4] <= fa_s0_c121_n944_c;
                    stage1_col122[5] <= fa_s0_c121_n945_c;
                    stage1_col122[6] <= fa_s0_c121_n946_c;
                    stage1_col122[7] <= fa_s0_c121_n947_c;
                    stage1_col122[8] <= fa_s0_c121_n948_c;
                    stage1_col122[9] <= fa_s0_c121_n949_c;
                    stage1_col122[10] <= fa_s0_c122_n950_s;
                    stage1_col122[11] <= fa_s0_c122_n951_s;
                    stage1_col122[12] <= fa_s0_c122_n952_s;
                    stage1_col122[13] <= fa_s0_c122_n953_s;
                    stage1_col122[14] <= fa_s0_c122_n954_s;
                    stage1_col122[15] <= fa_s0_c122_n955_s;
                    stage1_col122[16] <= fa_s0_c122_n956_s;
                    stage1_col122[17] <= fa_s0_c122_n957_s;
                    stage1_col122[18] <= fa_s0_c122_n958_s;
                    stage1_col122[19] <= fa_s0_c122_n959_s;
                    stage1_col122[20] <= fa_s0_c122_n960_s;
                    stage1_col123[0] <= fa_s0_c122_n950_c;
                    stage1_col123[1] <= fa_s0_c122_n951_c;
                    stage1_col123[2] <= fa_s0_c122_n952_c;
                    stage1_col123[3] <= fa_s0_c122_n953_c;
                    stage1_col123[4] <= fa_s0_c122_n954_c;
                    stage1_col123[5] <= fa_s0_c122_n955_c;
                    stage1_col123[6] <= fa_s0_c122_n956_c;
                    stage1_col123[7] <= fa_s0_c122_n957_c;
                    stage1_col123[8] <= fa_s0_c122_n958_c;
                    stage1_col123[9] <= fa_s0_c122_n959_c;
                    stage1_col123[10] <= fa_s0_c122_n960_c;
                    stage1_col123[11] <= fa_s0_c123_n961_s;
                    stage1_col123[12] <= fa_s0_c123_n962_s;
                    stage1_col123[13] <= fa_s0_c123_n963_s;
                    stage1_col123[14] <= fa_s0_c123_n964_s;
                    stage1_col123[15] <= fa_s0_c123_n965_s;
                    stage1_col123[16] <= fa_s0_c123_n966_s;
                    stage1_col123[17] <= fa_s0_c123_n967_s;
                    stage1_col123[18] <= fa_s0_c123_n968_s;
                    stage1_col123[19] <= fa_s0_c123_n969_s;
                    stage1_col123[20] <= fa_s0_c123_n970_s;
                    stage1_col123[21] <= stage0_col123[30];
                    stage1_col123[22] <= stage0_col123[31];
                    stage1_col124[0] <= fa_s0_c123_n961_c;
                    stage1_col124[1] <= fa_s0_c123_n962_c;
                    stage1_col124[2] <= fa_s0_c123_n963_c;
                    stage1_col124[3] <= fa_s0_c123_n964_c;
                    stage1_col124[4] <= fa_s0_c123_n965_c;
                    stage1_col124[5] <= fa_s0_c123_n966_c;
                    stage1_col124[6] <= fa_s0_c123_n967_c;
                    stage1_col124[7] <= fa_s0_c123_n968_c;
                    stage1_col124[8] <= fa_s0_c123_n969_c;
                    stage1_col124[9] <= fa_s0_c123_n970_c;
                    stage1_col124[10] <= fa_s0_c124_n971_s;
                    stage1_col124[11] <= fa_s0_c124_n972_s;
                    stage1_col124[12] <= fa_s0_c124_n973_s;
                    stage1_col124[13] <= fa_s0_c124_n974_s;
                    stage1_col124[14] <= fa_s0_c124_n975_s;
                    stage1_col124[15] <= fa_s0_c124_n976_s;
                    stage1_col124[16] <= fa_s0_c124_n977_s;
                    stage1_col124[17] <= fa_s0_c124_n978_s;
                    stage1_col124[18] <= fa_s0_c124_n979_s;
                    stage1_col124[19] <= fa_s0_c124_n980_s;
                    stage1_col124[20] <= fa_s0_c124_n981_s;
                    stage1_col125[0] <= fa_s0_c124_n971_c;
                    stage1_col125[1] <= fa_s0_c124_n972_c;
                    stage1_col125[2] <= fa_s0_c124_n973_c;
                    stage1_col125[3] <= fa_s0_c124_n974_c;
                    stage1_col125[4] <= fa_s0_c124_n975_c;
                    stage1_col125[5] <= fa_s0_c124_n976_c;
                    stage1_col125[6] <= fa_s0_c124_n977_c;
                    stage1_col125[7] <= fa_s0_c124_n978_c;
                    stage1_col125[8] <= fa_s0_c124_n979_c;
                    stage1_col125[9] <= fa_s0_c124_n980_c;
                    stage1_col125[10] <= fa_s0_c124_n981_c;
                    stage1_col125[11] <= fa_s0_c125_n982_s;
                    stage1_col125[12] <= fa_s0_c125_n983_s;
                    stage1_col125[13] <= fa_s0_c125_n984_s;
                    stage1_col125[14] <= fa_s0_c125_n985_s;
                    stage1_col125[15] <= fa_s0_c125_n986_s;
                    stage1_col125[16] <= fa_s0_c125_n987_s;
                    stage1_col125[17] <= fa_s0_c125_n988_s;
                    stage1_col125[18] <= fa_s0_c125_n989_s;
                    stage1_col125[19] <= fa_s0_c125_n990_s;
                    stage1_col125[20] <= fa_s0_c125_n991_s;
                    stage1_col125[21] <= stage0_col125[0];
                    stage1_col125[22] <= stage0_col125[31];
                    stage1_col126[0] <= fa_s0_c125_n982_c;
                    stage1_col126[1] <= fa_s0_c125_n983_c;
                    stage1_col126[2] <= fa_s0_c125_n984_c;
                    stage1_col126[3] <= fa_s0_c125_n985_c;
                    stage1_col126[4] <= fa_s0_c125_n986_c;
                    stage1_col126[5] <= fa_s0_c125_n987_c;
                    stage1_col126[6] <= fa_s0_c125_n988_c;
                    stage1_col126[7] <= fa_s0_c125_n989_c;
                    stage1_col126[8] <= fa_s0_c125_n990_c;
                    stage1_col126[9] <= fa_s0_c125_n991_c;
                    stage1_col126[10] <= fa_s0_c126_n992_s;
                    stage1_col126[11] <= fa_s0_c126_n993_s;
                    stage1_col126[12] <= fa_s0_c126_n994_s;
                    stage1_col126[13] <= fa_s0_c126_n995_s;
                    stage1_col126[14] <= fa_s0_c126_n996_s;
                    stage1_col126[15] <= fa_s0_c126_n997_s;
                    stage1_col126[16] <= fa_s0_c126_n998_s;
                    stage1_col126[17] <= fa_s0_c126_n999_s;
                    stage1_col126[18] <= fa_s0_c126_n1000_s;
                    stage1_col126[19] <= fa_s0_c126_n1001_s;
                    stage1_col126[20] <= fa_s0_c126_n1002_s;
                    stage1_col127[0] <= fa_s0_c126_n992_c;
                    stage1_col127[1] <= fa_s0_c126_n993_c;
                    stage1_col127[2] <= fa_s0_c126_n994_c;
                    stage1_col127[3] <= fa_s0_c126_n995_c;
                    stage1_col127[4] <= fa_s0_c126_n996_c;
                    stage1_col127[5] <= fa_s0_c126_n997_c;
                    stage1_col127[6] <= fa_s0_c126_n998_c;
                    stage1_col127[7] <= fa_s0_c126_n999_c;
                    stage1_col127[8] <= fa_s0_c126_n1000_c;
                    stage1_col127[9] <= fa_s0_c126_n1001_c;
                    stage1_col127[10] <= fa_s0_c126_n1002_c;
                    stage1_col127[11] <= stage0_col127[0];
                    stage1_col127[12] <= stage0_col127[0];
                    stage1_col127[13] <= stage0_col127[0];
                    stage1_col127[14] <= stage0_col127[0];
                    stage1_col127[15] <= stage0_col127[0];
                    stage1_col127[16] <= stage0_col127[0];
                    stage1_col127[17] <= stage0_col127[0];
                    stage1_col127[18] <= stage0_col127[0];
                    stage1_col127[19] <= stage0_col127[0];
                    stage1_col127[20] <= stage0_col127[0];
                    stage1_col127[21] <= stage0_col127[0];
                    stage1_col127[22] <= stage0_col127[0];
                    stage1_col127[23] <= stage0_col127[0];
                    stage1_col127[24] <= stage0_col127[0];
                    stage1_col127[25] <= stage0_col127[0];
                    stage1_col127[26] <= stage0_col127[0];
                    stage1_col127[27] <= stage0_col127[0];
                    stage1_col127[28] <= stage0_col127[0];
                    stage1_col127[29] <= stage0_col127[0];
                    stage1_col127[30] <= stage0_col127[0];
                    stage1_col127[31] <= stage0_col127[0];
                    stage1_col127[32] <= stage0_col127[0];
                    stage1_col127[33] <= stage0_col127[0];
                    stage1_col127[34] <= stage0_col127[0];
                    stage1_col127[35] <= stage0_col127[0];
                    stage1_col127[36] <= stage0_col127[0];
                    stage1_col127[37] <= stage0_col127[0];
                    stage1_col127[38] <= stage0_col127[0];
                    stage1_col127[39] <= stage0_col127[0];
                    stage1_col127[40] <= stage0_col127[0];
                    stage1_col127[41] <= stage0_col127[0];
                    stage1_col127[42] <= stage0_col127[0];
                end
            end
        end else begin : gen_stage1_no_pipe
            // Combinational assignment
            always_comb begin
                stage1_col0[0] = ha_s0_c0_n0_s;
                stage1_col1[0] = ha_s0_c0_n0_c;
                stage1_col1[1] = stage0_col1[0];
                stage1_col2[0] = fa_s0_c2_n0_s;
                stage1_col3[0] = fa_s0_c2_n0_c;
                stage1_col3[1] = stage0_col3[0];
                stage1_col3[2] = stage0_col3[1];
                stage1_col4[0] = fa_s0_c4_n1_s;
                stage1_col4[1] = stage0_col4[3];
                stage1_col5[0] = fa_s0_c4_n1_c;
                stage1_col5[1] = fa_s0_c5_n2_s;
                stage1_col6[0] = fa_s0_c5_n2_c;
                stage1_col6[1] = fa_s0_c6_n3_s;
                stage1_col6[2] = stage0_col6[3];
                stage1_col6[3] = stage0_col6[4];
                stage1_col7[0] = fa_s0_c6_n3_c;
                stage1_col7[1] = fa_s0_c7_n4_s;
                stage1_col7[2] = stage0_col7[3];
                stage1_col8[0] = fa_s0_c7_n4_c;
                stage1_col8[1] = fa_s0_c8_n5_s;
                stage1_col8[2] = fa_s0_c8_n6_s;
                stage1_col9[0] = fa_s0_c8_n5_c;
                stage1_col9[1] = fa_s0_c8_n6_c;
                stage1_col9[2] = fa_s0_c9_n7_s;
                stage1_col9[3] = stage0_col9[3];
                stage1_col9[4] = stage0_col9[4];
                stage1_col10[0] = fa_s0_c9_n7_c;
                stage1_col10[1] = fa_s0_c10_n8_s;
                stage1_col10[2] = fa_s0_c10_n9_s;
                stage1_col10[3] = stage0_col10[6];
                stage1_col11[0] = fa_s0_c10_n8_c;
                stage1_col11[1] = fa_s0_c10_n9_c;
                stage1_col11[2] = fa_s0_c11_n10_s;
                stage1_col11[3] = fa_s0_c11_n11_s;
                stage1_col12[0] = fa_s0_c11_n10_c;
                stage1_col12[1] = fa_s0_c11_n11_c;
                stage1_col12[2] = fa_s0_c12_n12_s;
                stage1_col12[3] = fa_s0_c12_n13_s;
                stage1_col12[4] = stage0_col12[6];
                stage1_col12[5] = stage0_col12[7];
                stage1_col13[0] = fa_s0_c12_n12_c;
                stage1_col13[1] = fa_s0_c12_n13_c;
                stage1_col13[2] = fa_s0_c13_n14_s;
                stage1_col13[3] = fa_s0_c13_n15_s;
                stage1_col13[4] = stage0_col13[6];
                stage1_col14[0] = fa_s0_c13_n14_c;
                stage1_col14[1] = fa_s0_c13_n15_c;
                stage1_col14[2] = fa_s0_c14_n16_s;
                stage1_col14[3] = fa_s0_c14_n17_s;
                stage1_col14[4] = fa_s0_c14_n18_s;
                stage1_col15[0] = fa_s0_c14_n16_c;
                stage1_col15[1] = fa_s0_c14_n17_c;
                stage1_col15[2] = fa_s0_c14_n18_c;
                stage1_col15[3] = fa_s0_c15_n19_s;
                stage1_col15[4] = fa_s0_c15_n20_s;
                stage1_col15[5] = stage0_col15[6];
                stage1_col15[6] = stage0_col15[7];
                stage1_col16[0] = fa_s0_c15_n19_c;
                stage1_col16[1] = fa_s0_c15_n20_c;
                stage1_col16[2] = fa_s0_c16_n21_s;
                stage1_col16[3] = fa_s0_c16_n22_s;
                stage1_col16[4] = fa_s0_c16_n23_s;
                stage1_col16[5] = stage0_col16[9];
                stage1_col17[0] = fa_s0_c16_n21_c;
                stage1_col17[1] = fa_s0_c16_n22_c;
                stage1_col17[2] = fa_s0_c16_n23_c;
                stage1_col17[3] = fa_s0_c17_n24_s;
                stage1_col17[4] = fa_s0_c17_n25_s;
                stage1_col17[5] = fa_s0_c17_n26_s;
                stage1_col18[0] = fa_s0_c17_n24_c;
                stage1_col18[1] = fa_s0_c17_n25_c;
                stage1_col18[2] = fa_s0_c17_n26_c;
                stage1_col18[3] = fa_s0_c18_n27_s;
                stage1_col18[4] = fa_s0_c18_n28_s;
                stage1_col18[5] = fa_s0_c18_n29_s;
                stage1_col18[6] = stage0_col18[9];
                stage1_col18[7] = stage0_col18[10];
                stage1_col19[0] = fa_s0_c18_n27_c;
                stage1_col19[1] = fa_s0_c18_n28_c;
                stage1_col19[2] = fa_s0_c18_n29_c;
                stage1_col19[3] = fa_s0_c19_n30_s;
                stage1_col19[4] = fa_s0_c19_n31_s;
                stage1_col19[5] = fa_s0_c19_n32_s;
                stage1_col19[6] = stage0_col19[9];
                stage1_col20[0] = fa_s0_c19_n30_c;
                stage1_col20[1] = fa_s0_c19_n31_c;
                stage1_col20[2] = fa_s0_c19_n32_c;
                stage1_col20[3] = fa_s0_c20_n33_s;
                stage1_col20[4] = fa_s0_c20_n34_s;
                stage1_col20[5] = fa_s0_c20_n35_s;
                stage1_col20[6] = fa_s0_c20_n36_s;
                stage1_col21[0] = fa_s0_c20_n33_c;
                stage1_col21[1] = fa_s0_c20_n34_c;
                stage1_col21[2] = fa_s0_c20_n35_c;
                stage1_col21[3] = fa_s0_c20_n36_c;
                stage1_col21[4] = fa_s0_c21_n37_s;
                stage1_col21[5] = fa_s0_c21_n38_s;
                stage1_col21[6] = fa_s0_c21_n39_s;
                stage1_col21[7] = stage0_col21[9];
                stage1_col21[8] = stage0_col21[10];
                stage1_col22[0] = fa_s0_c21_n37_c;
                stage1_col22[1] = fa_s0_c21_n38_c;
                stage1_col22[2] = fa_s0_c21_n39_c;
                stage1_col22[3] = fa_s0_c22_n40_s;
                stage1_col22[4] = fa_s0_c22_n41_s;
                stage1_col22[5] = fa_s0_c22_n42_s;
                stage1_col22[6] = fa_s0_c22_n43_s;
                stage1_col22[7] = stage0_col22[12];
                stage1_col23[0] = fa_s0_c22_n40_c;
                stage1_col23[1] = fa_s0_c22_n41_c;
                stage1_col23[2] = fa_s0_c22_n42_c;
                stage1_col23[3] = fa_s0_c22_n43_c;
                stage1_col23[4] = fa_s0_c23_n44_s;
                stage1_col23[5] = fa_s0_c23_n45_s;
                stage1_col23[6] = fa_s0_c23_n46_s;
                stage1_col23[7] = fa_s0_c23_n47_s;
                stage1_col24[0] = fa_s0_c23_n44_c;
                stage1_col24[1] = fa_s0_c23_n45_c;
                stage1_col24[2] = fa_s0_c23_n46_c;
                stage1_col24[3] = fa_s0_c23_n47_c;
                stage1_col24[4] = fa_s0_c24_n48_s;
                stage1_col24[5] = fa_s0_c24_n49_s;
                stage1_col24[6] = fa_s0_c24_n50_s;
                stage1_col24[7] = fa_s0_c24_n51_s;
                stage1_col24[8] = stage0_col24[12];
                stage1_col24[9] = stage0_col24[13];
                stage1_col25[0] = fa_s0_c24_n48_c;
                stage1_col25[1] = fa_s0_c24_n49_c;
                stage1_col25[2] = fa_s0_c24_n50_c;
                stage1_col25[3] = fa_s0_c24_n51_c;
                stage1_col25[4] = fa_s0_c25_n52_s;
                stage1_col25[5] = fa_s0_c25_n53_s;
                stage1_col25[6] = fa_s0_c25_n54_s;
                stage1_col25[7] = fa_s0_c25_n55_s;
                stage1_col25[8] = stage0_col25[12];
                stage1_col26[0] = fa_s0_c25_n52_c;
                stage1_col26[1] = fa_s0_c25_n53_c;
                stage1_col26[2] = fa_s0_c25_n54_c;
                stage1_col26[3] = fa_s0_c25_n55_c;
                stage1_col26[4] = fa_s0_c26_n56_s;
                stage1_col26[5] = fa_s0_c26_n57_s;
                stage1_col26[6] = fa_s0_c26_n58_s;
                stage1_col26[7] = fa_s0_c26_n59_s;
                stage1_col26[8] = fa_s0_c26_n60_s;
                stage1_col27[0] = fa_s0_c26_n56_c;
                stage1_col27[1] = fa_s0_c26_n57_c;
                stage1_col27[2] = fa_s0_c26_n58_c;
                stage1_col27[3] = fa_s0_c26_n59_c;
                stage1_col27[4] = fa_s0_c26_n60_c;
                stage1_col27[5] = fa_s0_c27_n61_s;
                stage1_col27[6] = fa_s0_c27_n62_s;
                stage1_col27[7] = fa_s0_c27_n63_s;
                stage1_col27[8] = fa_s0_c27_n64_s;
                stage1_col27[9] = stage0_col27[12];
                stage1_col27[10] = stage0_col27[13];
                stage1_col28[0] = fa_s0_c27_n61_c;
                stage1_col28[1] = fa_s0_c27_n62_c;
                stage1_col28[2] = fa_s0_c27_n63_c;
                stage1_col28[3] = fa_s0_c27_n64_c;
                stage1_col28[4] = fa_s0_c28_n65_s;
                stage1_col28[5] = fa_s0_c28_n66_s;
                stage1_col28[6] = fa_s0_c28_n67_s;
                stage1_col28[7] = fa_s0_c28_n68_s;
                stage1_col28[8] = fa_s0_c28_n69_s;
                stage1_col28[9] = stage0_col28[15];
                stage1_col29[0] = fa_s0_c28_n65_c;
                stage1_col29[1] = fa_s0_c28_n66_c;
                stage1_col29[2] = fa_s0_c28_n67_c;
                stage1_col29[3] = fa_s0_c28_n68_c;
                stage1_col29[4] = fa_s0_c28_n69_c;
                stage1_col29[5] = fa_s0_c29_n70_s;
                stage1_col29[6] = fa_s0_c29_n71_s;
                stage1_col29[7] = fa_s0_c29_n72_s;
                stage1_col29[8] = fa_s0_c29_n73_s;
                stage1_col29[9] = fa_s0_c29_n74_s;
                stage1_col30[0] = fa_s0_c29_n70_c;
                stage1_col30[1] = fa_s0_c29_n71_c;
                stage1_col30[2] = fa_s0_c29_n72_c;
                stage1_col30[3] = fa_s0_c29_n73_c;
                stage1_col30[4] = fa_s0_c29_n74_c;
                stage1_col30[5] = fa_s0_c30_n75_s;
                stage1_col30[6] = fa_s0_c30_n76_s;
                stage1_col30[7] = fa_s0_c30_n77_s;
                stage1_col30[8] = fa_s0_c30_n78_s;
                stage1_col30[9] = fa_s0_c30_n79_s;
                stage1_col30[10] = stage0_col30[15];
                stage1_col30[11] = stage0_col30[16];
                stage1_col31[0] = fa_s0_c30_n75_c;
                stage1_col31[1] = fa_s0_c30_n76_c;
                stage1_col31[2] = fa_s0_c30_n77_c;
                stage1_col31[3] = fa_s0_c30_n78_c;
                stage1_col31[4] = fa_s0_c30_n79_c;
                stage1_col31[5] = fa_s0_c31_n80_s;
                stage1_col31[6] = fa_s0_c31_n81_s;
                stage1_col31[7] = fa_s0_c31_n82_s;
                stage1_col31[8] = fa_s0_c31_n83_s;
                stage1_col31[9] = fa_s0_c31_n84_s;
                stage1_col31[10] = stage0_col31[15];
                stage1_col32[0] = fa_s0_c31_n80_c;
                stage1_col32[1] = fa_s0_c31_n81_c;
                stage1_col32[2] = fa_s0_c31_n82_c;
                stage1_col32[3] = fa_s0_c31_n83_c;
                stage1_col32[4] = fa_s0_c31_n84_c;
                stage1_col32[5] = fa_s0_c32_n85_s;
                stage1_col32[6] = fa_s0_c32_n86_s;
                stage1_col32[7] = fa_s0_c32_n87_s;
                stage1_col32[8] = fa_s0_c32_n88_s;
                stage1_col32[9] = fa_s0_c32_n89_s;
                stage1_col32[10] = fa_s0_c32_n90_s;
                stage1_col33[0] = fa_s0_c32_n85_c;
                stage1_col33[1] = fa_s0_c32_n86_c;
                stage1_col33[2] = fa_s0_c32_n87_c;
                stage1_col33[3] = fa_s0_c32_n88_c;
                stage1_col33[4] = fa_s0_c32_n89_c;
                stage1_col33[5] = fa_s0_c32_n90_c;
                stage1_col33[6] = fa_s0_c33_n91_s;
                stage1_col33[7] = fa_s0_c33_n92_s;
                stage1_col33[8] = fa_s0_c33_n93_s;
                stage1_col33[9] = fa_s0_c33_n94_s;
                stage1_col33[10] = fa_s0_c33_n95_s;
                stage1_col33[11] = stage0_col33[15];
                stage1_col33[12] = stage0_col33[16];
                stage1_col34[0] = fa_s0_c33_n91_c;
                stage1_col34[1] = fa_s0_c33_n92_c;
                stage1_col34[2] = fa_s0_c33_n93_c;
                stage1_col34[3] = fa_s0_c33_n94_c;
                stage1_col34[4] = fa_s0_c33_n95_c;
                stage1_col34[5] = fa_s0_c34_n96_s;
                stage1_col34[6] = fa_s0_c34_n97_s;
                stage1_col34[7] = fa_s0_c34_n98_s;
                stage1_col34[8] = fa_s0_c34_n99_s;
                stage1_col34[9] = fa_s0_c34_n100_s;
                stage1_col34[10] = fa_s0_c34_n101_s;
                stage1_col34[11] = stage0_col34[18];
                stage1_col35[0] = fa_s0_c34_n96_c;
                stage1_col35[1] = fa_s0_c34_n97_c;
                stage1_col35[2] = fa_s0_c34_n98_c;
                stage1_col35[3] = fa_s0_c34_n99_c;
                stage1_col35[4] = fa_s0_c34_n100_c;
                stage1_col35[5] = fa_s0_c34_n101_c;
                stage1_col35[6] = fa_s0_c35_n102_s;
                stage1_col35[7] = fa_s0_c35_n103_s;
                stage1_col35[8] = fa_s0_c35_n104_s;
                stage1_col35[9] = fa_s0_c35_n105_s;
                stage1_col35[10] = fa_s0_c35_n106_s;
                stage1_col35[11] = fa_s0_c35_n107_s;
                stage1_col36[0] = fa_s0_c35_n102_c;
                stage1_col36[1] = fa_s0_c35_n103_c;
                stage1_col36[2] = fa_s0_c35_n104_c;
                stage1_col36[3] = fa_s0_c35_n105_c;
                stage1_col36[4] = fa_s0_c35_n106_c;
                stage1_col36[5] = fa_s0_c35_n107_c;
                stage1_col36[6] = fa_s0_c36_n108_s;
                stage1_col36[7] = fa_s0_c36_n109_s;
                stage1_col36[8] = fa_s0_c36_n110_s;
                stage1_col36[9] = fa_s0_c36_n111_s;
                stage1_col36[10] = fa_s0_c36_n112_s;
                stage1_col36[11] = fa_s0_c36_n113_s;
                stage1_col36[12] = stage0_col36[18];
                stage1_col36[13] = stage0_col36[19];
                stage1_col37[0] = fa_s0_c36_n108_c;
                stage1_col37[1] = fa_s0_c36_n109_c;
                stage1_col37[2] = fa_s0_c36_n110_c;
                stage1_col37[3] = fa_s0_c36_n111_c;
                stage1_col37[4] = fa_s0_c36_n112_c;
                stage1_col37[5] = fa_s0_c36_n113_c;
                stage1_col37[6] = fa_s0_c37_n114_s;
                stage1_col37[7] = fa_s0_c37_n115_s;
                stage1_col37[8] = fa_s0_c37_n116_s;
                stage1_col37[9] = fa_s0_c37_n117_s;
                stage1_col37[10] = fa_s0_c37_n118_s;
                stage1_col37[11] = fa_s0_c37_n119_s;
                stage1_col37[12] = stage0_col37[18];
                stage1_col38[0] = fa_s0_c37_n114_c;
                stage1_col38[1] = fa_s0_c37_n115_c;
                stage1_col38[2] = fa_s0_c37_n116_c;
                stage1_col38[3] = fa_s0_c37_n117_c;
                stage1_col38[4] = fa_s0_c37_n118_c;
                stage1_col38[5] = fa_s0_c37_n119_c;
                stage1_col38[6] = fa_s0_c38_n120_s;
                stage1_col38[7] = fa_s0_c38_n121_s;
                stage1_col38[8] = fa_s0_c38_n122_s;
                stage1_col38[9] = fa_s0_c38_n123_s;
                stage1_col38[10] = fa_s0_c38_n124_s;
                stage1_col38[11] = fa_s0_c38_n125_s;
                stage1_col38[12] = fa_s0_c38_n126_s;
                stage1_col39[0] = fa_s0_c38_n120_c;
                stage1_col39[1] = fa_s0_c38_n121_c;
                stage1_col39[2] = fa_s0_c38_n122_c;
                stage1_col39[3] = fa_s0_c38_n123_c;
                stage1_col39[4] = fa_s0_c38_n124_c;
                stage1_col39[5] = fa_s0_c38_n125_c;
                stage1_col39[6] = fa_s0_c38_n126_c;
                stage1_col39[7] = fa_s0_c39_n127_s;
                stage1_col39[8] = fa_s0_c39_n128_s;
                stage1_col39[9] = fa_s0_c39_n129_s;
                stage1_col39[10] = fa_s0_c39_n130_s;
                stage1_col39[11] = fa_s0_c39_n131_s;
                stage1_col39[12] = fa_s0_c39_n132_s;
                stage1_col39[13] = stage0_col39[18];
                stage1_col39[14] = stage0_col39[19];
                stage1_col40[0] = fa_s0_c39_n127_c;
                stage1_col40[1] = fa_s0_c39_n128_c;
                stage1_col40[2] = fa_s0_c39_n129_c;
                stage1_col40[3] = fa_s0_c39_n130_c;
                stage1_col40[4] = fa_s0_c39_n131_c;
                stage1_col40[5] = fa_s0_c39_n132_c;
                stage1_col40[6] = fa_s0_c40_n133_s;
                stage1_col40[7] = fa_s0_c40_n134_s;
                stage1_col40[8] = fa_s0_c40_n135_s;
                stage1_col40[9] = fa_s0_c40_n136_s;
                stage1_col40[10] = fa_s0_c40_n137_s;
                stage1_col40[11] = fa_s0_c40_n138_s;
                stage1_col40[12] = fa_s0_c40_n139_s;
                stage1_col40[13] = stage0_col40[21];
                stage1_col41[0] = fa_s0_c40_n133_c;
                stage1_col41[1] = fa_s0_c40_n134_c;
                stage1_col41[2] = fa_s0_c40_n135_c;
                stage1_col41[3] = fa_s0_c40_n136_c;
                stage1_col41[4] = fa_s0_c40_n137_c;
                stage1_col41[5] = fa_s0_c40_n138_c;
                stage1_col41[6] = fa_s0_c40_n139_c;
                stage1_col41[7] = fa_s0_c41_n140_s;
                stage1_col41[8] = fa_s0_c41_n141_s;
                stage1_col41[9] = fa_s0_c41_n142_s;
                stage1_col41[10] = fa_s0_c41_n143_s;
                stage1_col41[11] = fa_s0_c41_n144_s;
                stage1_col41[12] = fa_s0_c41_n145_s;
                stage1_col41[13] = fa_s0_c41_n146_s;
                stage1_col42[0] = fa_s0_c41_n140_c;
                stage1_col42[1] = fa_s0_c41_n141_c;
                stage1_col42[2] = fa_s0_c41_n142_c;
                stage1_col42[3] = fa_s0_c41_n143_c;
                stage1_col42[4] = fa_s0_c41_n144_c;
                stage1_col42[5] = fa_s0_c41_n145_c;
                stage1_col42[6] = fa_s0_c41_n146_c;
                stage1_col42[7] = fa_s0_c42_n147_s;
                stage1_col42[8] = fa_s0_c42_n148_s;
                stage1_col42[9] = fa_s0_c42_n149_s;
                stage1_col42[10] = fa_s0_c42_n150_s;
                stage1_col42[11] = fa_s0_c42_n151_s;
                stage1_col42[12] = fa_s0_c42_n152_s;
                stage1_col42[13] = fa_s0_c42_n153_s;
                stage1_col42[14] = stage0_col42[21];
                stage1_col42[15] = stage0_col42[22];
                stage1_col43[0] = fa_s0_c42_n147_c;
                stage1_col43[1] = fa_s0_c42_n148_c;
                stage1_col43[2] = fa_s0_c42_n149_c;
                stage1_col43[3] = fa_s0_c42_n150_c;
                stage1_col43[4] = fa_s0_c42_n151_c;
                stage1_col43[5] = fa_s0_c42_n152_c;
                stage1_col43[6] = fa_s0_c42_n153_c;
                stage1_col43[7] = fa_s0_c43_n154_s;
                stage1_col43[8] = fa_s0_c43_n155_s;
                stage1_col43[9] = fa_s0_c43_n156_s;
                stage1_col43[10] = fa_s0_c43_n157_s;
                stage1_col43[11] = fa_s0_c43_n158_s;
                stage1_col43[12] = fa_s0_c43_n159_s;
                stage1_col43[13] = fa_s0_c43_n160_s;
                stage1_col43[14] = stage0_col43[21];
                stage1_col44[0] = fa_s0_c43_n154_c;
                stage1_col44[1] = fa_s0_c43_n155_c;
                stage1_col44[2] = fa_s0_c43_n156_c;
                stage1_col44[3] = fa_s0_c43_n157_c;
                stage1_col44[4] = fa_s0_c43_n158_c;
                stage1_col44[5] = fa_s0_c43_n159_c;
                stage1_col44[6] = fa_s0_c43_n160_c;
                stage1_col44[7] = fa_s0_c44_n161_s;
                stage1_col44[8] = fa_s0_c44_n162_s;
                stage1_col44[9] = fa_s0_c44_n163_s;
                stage1_col44[10] = fa_s0_c44_n164_s;
                stage1_col44[11] = fa_s0_c44_n165_s;
                stage1_col44[12] = fa_s0_c44_n166_s;
                stage1_col44[13] = fa_s0_c44_n167_s;
                stage1_col44[14] = fa_s0_c44_n168_s;
                stage1_col45[0] = fa_s0_c44_n161_c;
                stage1_col45[1] = fa_s0_c44_n162_c;
                stage1_col45[2] = fa_s0_c44_n163_c;
                stage1_col45[3] = fa_s0_c44_n164_c;
                stage1_col45[4] = fa_s0_c44_n165_c;
                stage1_col45[5] = fa_s0_c44_n166_c;
                stage1_col45[6] = fa_s0_c44_n167_c;
                stage1_col45[7] = fa_s0_c44_n168_c;
                stage1_col45[8] = fa_s0_c45_n169_s;
                stage1_col45[9] = fa_s0_c45_n170_s;
                stage1_col45[10] = fa_s0_c45_n171_s;
                stage1_col45[11] = fa_s0_c45_n172_s;
                stage1_col45[12] = fa_s0_c45_n173_s;
                stage1_col45[13] = fa_s0_c45_n174_s;
                stage1_col45[14] = fa_s0_c45_n175_s;
                stage1_col45[15] = stage0_col45[21];
                stage1_col45[16] = stage0_col45[22];
                stage1_col46[0] = fa_s0_c45_n169_c;
                stage1_col46[1] = fa_s0_c45_n170_c;
                stage1_col46[2] = fa_s0_c45_n171_c;
                stage1_col46[3] = fa_s0_c45_n172_c;
                stage1_col46[4] = fa_s0_c45_n173_c;
                stage1_col46[5] = fa_s0_c45_n174_c;
                stage1_col46[6] = fa_s0_c45_n175_c;
                stage1_col46[7] = fa_s0_c46_n176_s;
                stage1_col46[8] = fa_s0_c46_n177_s;
                stage1_col46[9] = fa_s0_c46_n178_s;
                stage1_col46[10] = fa_s0_c46_n179_s;
                stage1_col46[11] = fa_s0_c46_n180_s;
                stage1_col46[12] = fa_s0_c46_n181_s;
                stage1_col46[13] = fa_s0_c46_n182_s;
                stage1_col46[14] = fa_s0_c46_n183_s;
                stage1_col46[15] = stage0_col46[24];
                stage1_col47[0] = fa_s0_c46_n176_c;
                stage1_col47[1] = fa_s0_c46_n177_c;
                stage1_col47[2] = fa_s0_c46_n178_c;
                stage1_col47[3] = fa_s0_c46_n179_c;
                stage1_col47[4] = fa_s0_c46_n180_c;
                stage1_col47[5] = fa_s0_c46_n181_c;
                stage1_col47[6] = fa_s0_c46_n182_c;
                stage1_col47[7] = fa_s0_c46_n183_c;
                stage1_col47[8] = fa_s0_c47_n184_s;
                stage1_col47[9] = fa_s0_c47_n185_s;
                stage1_col47[10] = fa_s0_c47_n186_s;
                stage1_col47[11] = fa_s0_c47_n187_s;
                stage1_col47[12] = fa_s0_c47_n188_s;
                stage1_col47[13] = fa_s0_c47_n189_s;
                stage1_col47[14] = fa_s0_c47_n190_s;
                stage1_col47[15] = fa_s0_c47_n191_s;
                stage1_col48[0] = fa_s0_c47_n184_c;
                stage1_col48[1] = fa_s0_c47_n185_c;
                stage1_col48[2] = fa_s0_c47_n186_c;
                stage1_col48[3] = fa_s0_c47_n187_c;
                stage1_col48[4] = fa_s0_c47_n188_c;
                stage1_col48[5] = fa_s0_c47_n189_c;
                stage1_col48[6] = fa_s0_c47_n190_c;
                stage1_col48[7] = fa_s0_c47_n191_c;
                stage1_col48[8] = fa_s0_c48_n192_s;
                stage1_col48[9] = fa_s0_c48_n193_s;
                stage1_col48[10] = fa_s0_c48_n194_s;
                stage1_col48[11] = fa_s0_c48_n195_s;
                stage1_col48[12] = fa_s0_c48_n196_s;
                stage1_col48[13] = fa_s0_c48_n197_s;
                stage1_col48[14] = fa_s0_c48_n198_s;
                stage1_col48[15] = fa_s0_c48_n199_s;
                stage1_col48[16] = stage0_col48[24];
                stage1_col48[17] = stage0_col48[25];
                stage1_col49[0] = fa_s0_c48_n192_c;
                stage1_col49[1] = fa_s0_c48_n193_c;
                stage1_col49[2] = fa_s0_c48_n194_c;
                stage1_col49[3] = fa_s0_c48_n195_c;
                stage1_col49[4] = fa_s0_c48_n196_c;
                stage1_col49[5] = fa_s0_c48_n197_c;
                stage1_col49[6] = fa_s0_c48_n198_c;
                stage1_col49[7] = fa_s0_c48_n199_c;
                stage1_col49[8] = fa_s0_c49_n200_s;
                stage1_col49[9] = fa_s0_c49_n201_s;
                stage1_col49[10] = fa_s0_c49_n202_s;
                stage1_col49[11] = fa_s0_c49_n203_s;
                stage1_col49[12] = fa_s0_c49_n204_s;
                stage1_col49[13] = fa_s0_c49_n205_s;
                stage1_col49[14] = fa_s0_c49_n206_s;
                stage1_col49[15] = fa_s0_c49_n207_s;
                stage1_col49[16] = stage0_col49[24];
                stage1_col50[0] = fa_s0_c49_n200_c;
                stage1_col50[1] = fa_s0_c49_n201_c;
                stage1_col50[2] = fa_s0_c49_n202_c;
                stage1_col50[3] = fa_s0_c49_n203_c;
                stage1_col50[4] = fa_s0_c49_n204_c;
                stage1_col50[5] = fa_s0_c49_n205_c;
                stage1_col50[6] = fa_s0_c49_n206_c;
                stage1_col50[7] = fa_s0_c49_n207_c;
                stage1_col50[8] = fa_s0_c50_n208_s;
                stage1_col50[9] = fa_s0_c50_n209_s;
                stage1_col50[10] = fa_s0_c50_n210_s;
                stage1_col50[11] = fa_s0_c50_n211_s;
                stage1_col50[12] = fa_s0_c50_n212_s;
                stage1_col50[13] = fa_s0_c50_n213_s;
                stage1_col50[14] = fa_s0_c50_n214_s;
                stage1_col50[15] = fa_s0_c50_n215_s;
                stage1_col50[16] = fa_s0_c50_n216_s;
                stage1_col51[0] = fa_s0_c50_n208_c;
                stage1_col51[1] = fa_s0_c50_n209_c;
                stage1_col51[2] = fa_s0_c50_n210_c;
                stage1_col51[3] = fa_s0_c50_n211_c;
                stage1_col51[4] = fa_s0_c50_n212_c;
                stage1_col51[5] = fa_s0_c50_n213_c;
                stage1_col51[6] = fa_s0_c50_n214_c;
                stage1_col51[7] = fa_s0_c50_n215_c;
                stage1_col51[8] = fa_s0_c50_n216_c;
                stage1_col51[9] = fa_s0_c51_n217_s;
                stage1_col51[10] = fa_s0_c51_n218_s;
                stage1_col51[11] = fa_s0_c51_n219_s;
                stage1_col51[12] = fa_s0_c51_n220_s;
                stage1_col51[13] = fa_s0_c51_n221_s;
                stage1_col51[14] = fa_s0_c51_n222_s;
                stage1_col51[15] = fa_s0_c51_n223_s;
                stage1_col51[16] = fa_s0_c51_n224_s;
                stage1_col51[17] = stage0_col51[24];
                stage1_col51[18] = stage0_col51[25];
                stage1_col52[0] = fa_s0_c51_n217_c;
                stage1_col52[1] = fa_s0_c51_n218_c;
                stage1_col52[2] = fa_s0_c51_n219_c;
                stage1_col52[3] = fa_s0_c51_n220_c;
                stage1_col52[4] = fa_s0_c51_n221_c;
                stage1_col52[5] = fa_s0_c51_n222_c;
                stage1_col52[6] = fa_s0_c51_n223_c;
                stage1_col52[7] = fa_s0_c51_n224_c;
                stage1_col52[8] = fa_s0_c52_n225_s;
                stage1_col52[9] = fa_s0_c52_n226_s;
                stage1_col52[10] = fa_s0_c52_n227_s;
                stage1_col52[11] = fa_s0_c52_n228_s;
                stage1_col52[12] = fa_s0_c52_n229_s;
                stage1_col52[13] = fa_s0_c52_n230_s;
                stage1_col52[14] = fa_s0_c52_n231_s;
                stage1_col52[15] = fa_s0_c52_n232_s;
                stage1_col52[16] = fa_s0_c52_n233_s;
                stage1_col52[17] = stage0_col52[27];
                stage1_col53[0] = fa_s0_c52_n225_c;
                stage1_col53[1] = fa_s0_c52_n226_c;
                stage1_col53[2] = fa_s0_c52_n227_c;
                stage1_col53[3] = fa_s0_c52_n228_c;
                stage1_col53[4] = fa_s0_c52_n229_c;
                stage1_col53[5] = fa_s0_c52_n230_c;
                stage1_col53[6] = fa_s0_c52_n231_c;
                stage1_col53[7] = fa_s0_c52_n232_c;
                stage1_col53[8] = fa_s0_c52_n233_c;
                stage1_col53[9] = fa_s0_c53_n234_s;
                stage1_col53[10] = fa_s0_c53_n235_s;
                stage1_col53[11] = fa_s0_c53_n236_s;
                stage1_col53[12] = fa_s0_c53_n237_s;
                stage1_col53[13] = fa_s0_c53_n238_s;
                stage1_col53[14] = fa_s0_c53_n239_s;
                stage1_col53[15] = fa_s0_c53_n240_s;
                stage1_col53[16] = fa_s0_c53_n241_s;
                stage1_col53[17] = fa_s0_c53_n242_s;
                stage1_col54[0] = fa_s0_c53_n234_c;
                stage1_col54[1] = fa_s0_c53_n235_c;
                stage1_col54[2] = fa_s0_c53_n236_c;
                stage1_col54[3] = fa_s0_c53_n237_c;
                stage1_col54[4] = fa_s0_c53_n238_c;
                stage1_col54[5] = fa_s0_c53_n239_c;
                stage1_col54[6] = fa_s0_c53_n240_c;
                stage1_col54[7] = fa_s0_c53_n241_c;
                stage1_col54[8] = fa_s0_c53_n242_c;
                stage1_col54[9] = fa_s0_c54_n243_s;
                stage1_col54[10] = fa_s0_c54_n244_s;
                stage1_col54[11] = fa_s0_c54_n245_s;
                stage1_col54[12] = fa_s0_c54_n246_s;
                stage1_col54[13] = fa_s0_c54_n247_s;
                stage1_col54[14] = fa_s0_c54_n248_s;
                stage1_col54[15] = fa_s0_c54_n249_s;
                stage1_col54[16] = fa_s0_c54_n250_s;
                stage1_col54[17] = fa_s0_c54_n251_s;
                stage1_col54[18] = stage0_col54[27];
                stage1_col54[19] = stage0_col54[28];
                stage1_col55[0] = fa_s0_c54_n243_c;
                stage1_col55[1] = fa_s0_c54_n244_c;
                stage1_col55[2] = fa_s0_c54_n245_c;
                stage1_col55[3] = fa_s0_c54_n246_c;
                stage1_col55[4] = fa_s0_c54_n247_c;
                stage1_col55[5] = fa_s0_c54_n248_c;
                stage1_col55[6] = fa_s0_c54_n249_c;
                stage1_col55[7] = fa_s0_c54_n250_c;
                stage1_col55[8] = fa_s0_c54_n251_c;
                stage1_col55[9] = fa_s0_c55_n252_s;
                stage1_col55[10] = fa_s0_c55_n253_s;
                stage1_col55[11] = fa_s0_c55_n254_s;
                stage1_col55[12] = fa_s0_c55_n255_s;
                stage1_col55[13] = fa_s0_c55_n256_s;
                stage1_col55[14] = fa_s0_c55_n257_s;
                stage1_col55[15] = fa_s0_c55_n258_s;
                stage1_col55[16] = fa_s0_c55_n259_s;
                stage1_col55[17] = fa_s0_c55_n260_s;
                stage1_col55[18] = stage0_col55[27];
                stage1_col56[0] = fa_s0_c55_n252_c;
                stage1_col56[1] = fa_s0_c55_n253_c;
                stage1_col56[2] = fa_s0_c55_n254_c;
                stage1_col56[3] = fa_s0_c55_n255_c;
                stage1_col56[4] = fa_s0_c55_n256_c;
                stage1_col56[5] = fa_s0_c55_n257_c;
                stage1_col56[6] = fa_s0_c55_n258_c;
                stage1_col56[7] = fa_s0_c55_n259_c;
                stage1_col56[8] = fa_s0_c55_n260_c;
                stage1_col56[9] = fa_s0_c56_n261_s;
                stage1_col56[10] = fa_s0_c56_n262_s;
                stage1_col56[11] = fa_s0_c56_n263_s;
                stage1_col56[12] = fa_s0_c56_n264_s;
                stage1_col56[13] = fa_s0_c56_n265_s;
                stage1_col56[14] = fa_s0_c56_n266_s;
                stage1_col56[15] = fa_s0_c56_n267_s;
                stage1_col56[16] = fa_s0_c56_n268_s;
                stage1_col56[17] = fa_s0_c56_n269_s;
                stage1_col56[18] = fa_s0_c56_n270_s;
                stage1_col57[0] = fa_s0_c56_n261_c;
                stage1_col57[1] = fa_s0_c56_n262_c;
                stage1_col57[2] = fa_s0_c56_n263_c;
                stage1_col57[3] = fa_s0_c56_n264_c;
                stage1_col57[4] = fa_s0_c56_n265_c;
                stage1_col57[5] = fa_s0_c56_n266_c;
                stage1_col57[6] = fa_s0_c56_n267_c;
                stage1_col57[7] = fa_s0_c56_n268_c;
                stage1_col57[8] = fa_s0_c56_n269_c;
                stage1_col57[9] = fa_s0_c56_n270_c;
                stage1_col57[10] = fa_s0_c57_n271_s;
                stage1_col57[11] = fa_s0_c57_n272_s;
                stage1_col57[12] = fa_s0_c57_n273_s;
                stage1_col57[13] = fa_s0_c57_n274_s;
                stage1_col57[14] = fa_s0_c57_n275_s;
                stage1_col57[15] = fa_s0_c57_n276_s;
                stage1_col57[16] = fa_s0_c57_n277_s;
                stage1_col57[17] = fa_s0_c57_n278_s;
                stage1_col57[18] = fa_s0_c57_n279_s;
                stage1_col57[19] = stage0_col57[27];
                stage1_col57[20] = stage0_col57[28];
                stage1_col58[0] = fa_s0_c57_n271_c;
                stage1_col58[1] = fa_s0_c57_n272_c;
                stage1_col58[2] = fa_s0_c57_n273_c;
                stage1_col58[3] = fa_s0_c57_n274_c;
                stage1_col58[4] = fa_s0_c57_n275_c;
                stage1_col58[5] = fa_s0_c57_n276_c;
                stage1_col58[6] = fa_s0_c57_n277_c;
                stage1_col58[7] = fa_s0_c57_n278_c;
                stage1_col58[8] = fa_s0_c57_n279_c;
                stage1_col58[9] = fa_s0_c58_n280_s;
                stage1_col58[10] = fa_s0_c58_n281_s;
                stage1_col58[11] = fa_s0_c58_n282_s;
                stage1_col58[12] = fa_s0_c58_n283_s;
                stage1_col58[13] = fa_s0_c58_n284_s;
                stage1_col58[14] = fa_s0_c58_n285_s;
                stage1_col58[15] = fa_s0_c58_n286_s;
                stage1_col58[16] = fa_s0_c58_n287_s;
                stage1_col58[17] = fa_s0_c58_n288_s;
                stage1_col58[18] = fa_s0_c58_n289_s;
                stage1_col58[19] = stage0_col58[30];
                stage1_col59[0] = fa_s0_c58_n280_c;
                stage1_col59[1] = fa_s0_c58_n281_c;
                stage1_col59[2] = fa_s0_c58_n282_c;
                stage1_col59[3] = fa_s0_c58_n283_c;
                stage1_col59[4] = fa_s0_c58_n284_c;
                stage1_col59[5] = fa_s0_c58_n285_c;
                stage1_col59[6] = fa_s0_c58_n286_c;
                stage1_col59[7] = fa_s0_c58_n287_c;
                stage1_col59[8] = fa_s0_c58_n288_c;
                stage1_col59[9] = fa_s0_c58_n289_c;
                stage1_col59[10] = fa_s0_c59_n290_s;
                stage1_col59[11] = fa_s0_c59_n291_s;
                stage1_col59[12] = fa_s0_c59_n292_s;
                stage1_col59[13] = fa_s0_c59_n293_s;
                stage1_col59[14] = fa_s0_c59_n294_s;
                stage1_col59[15] = fa_s0_c59_n295_s;
                stage1_col59[16] = fa_s0_c59_n296_s;
                stage1_col59[17] = fa_s0_c59_n297_s;
                stage1_col59[18] = fa_s0_c59_n298_s;
                stage1_col59[19] = fa_s0_c59_n299_s;
                stage1_col60[0] = fa_s0_c59_n290_c;
                stage1_col60[1] = fa_s0_c59_n291_c;
                stage1_col60[2] = fa_s0_c59_n292_c;
                stage1_col60[3] = fa_s0_c59_n293_c;
                stage1_col60[4] = fa_s0_c59_n294_c;
                stage1_col60[5] = fa_s0_c59_n295_c;
                stage1_col60[6] = fa_s0_c59_n296_c;
                stage1_col60[7] = fa_s0_c59_n297_c;
                stage1_col60[8] = fa_s0_c59_n298_c;
                stage1_col60[9] = fa_s0_c59_n299_c;
                stage1_col60[10] = fa_s0_c60_n300_s;
                stage1_col60[11] = fa_s0_c60_n301_s;
                stage1_col60[12] = fa_s0_c60_n302_s;
                stage1_col60[13] = fa_s0_c60_n303_s;
                stage1_col60[14] = fa_s0_c60_n304_s;
                stage1_col60[15] = fa_s0_c60_n305_s;
                stage1_col60[16] = fa_s0_c60_n306_s;
                stage1_col60[17] = fa_s0_c60_n307_s;
                stage1_col60[18] = fa_s0_c60_n308_s;
                stage1_col60[19] = fa_s0_c60_n309_s;
                stage1_col60[20] = stage0_col60[30];
                stage1_col60[21] = stage0_col60[31];
                stage1_col61[0] = fa_s0_c60_n300_c;
                stage1_col61[1] = fa_s0_c60_n301_c;
                stage1_col61[2] = fa_s0_c60_n302_c;
                stage1_col61[3] = fa_s0_c60_n303_c;
                stage1_col61[4] = fa_s0_c60_n304_c;
                stage1_col61[5] = fa_s0_c60_n305_c;
                stage1_col61[6] = fa_s0_c60_n306_c;
                stage1_col61[7] = fa_s0_c60_n307_c;
                stage1_col61[8] = fa_s0_c60_n308_c;
                stage1_col61[9] = fa_s0_c60_n309_c;
                stage1_col61[10] = fa_s0_c61_n310_s;
                stage1_col61[11] = fa_s0_c61_n311_s;
                stage1_col61[12] = fa_s0_c61_n312_s;
                stage1_col61[13] = fa_s0_c61_n313_s;
                stage1_col61[14] = fa_s0_c61_n314_s;
                stage1_col61[15] = fa_s0_c61_n315_s;
                stage1_col61[16] = fa_s0_c61_n316_s;
                stage1_col61[17] = fa_s0_c61_n317_s;
                stage1_col61[18] = fa_s0_c61_n318_s;
                stage1_col61[19] = fa_s0_c61_n319_s;
                stage1_col61[20] = stage0_col61[30];
                stage1_col62[0] = fa_s0_c61_n310_c;
                stage1_col62[1] = fa_s0_c61_n311_c;
                stage1_col62[2] = fa_s0_c61_n312_c;
                stage1_col62[3] = fa_s0_c61_n313_c;
                stage1_col62[4] = fa_s0_c61_n314_c;
                stage1_col62[5] = fa_s0_c61_n315_c;
                stage1_col62[6] = fa_s0_c61_n316_c;
                stage1_col62[7] = fa_s0_c61_n317_c;
                stage1_col62[8] = fa_s0_c61_n318_c;
                stage1_col62[9] = fa_s0_c61_n319_c;
                stage1_col62[10] = fa_s0_c62_n320_s;
                stage1_col62[11] = fa_s0_c62_n321_s;
                stage1_col62[12] = fa_s0_c62_n322_s;
                stage1_col62[13] = fa_s0_c62_n323_s;
                stage1_col62[14] = fa_s0_c62_n324_s;
                stage1_col62[15] = fa_s0_c62_n325_s;
                stage1_col62[16] = fa_s0_c62_n326_s;
                stage1_col62[17] = fa_s0_c62_n327_s;
                stage1_col62[18] = fa_s0_c62_n328_s;
                stage1_col62[19] = fa_s0_c62_n329_s;
                stage1_col62[20] = fa_s0_c62_n330_s;
                stage1_col63[0] = fa_s0_c62_n320_c;
                stage1_col63[1] = fa_s0_c62_n321_c;
                stage1_col63[2] = fa_s0_c62_n322_c;
                stage1_col63[3] = fa_s0_c62_n323_c;
                stage1_col63[4] = fa_s0_c62_n324_c;
                stage1_col63[5] = fa_s0_c62_n325_c;
                stage1_col63[6] = fa_s0_c62_n326_c;
                stage1_col63[7] = fa_s0_c62_n327_c;
                stage1_col63[8] = fa_s0_c62_n328_c;
                stage1_col63[9] = fa_s0_c62_n329_c;
                stage1_col63[10] = fa_s0_c62_n330_c;
                stage1_col63[11] = fa_s0_c63_n331_s;
                stage1_col63[12] = fa_s0_c63_n332_s;
                stage1_col63[13] = fa_s0_c63_n333_s;
                stage1_col63[14] = fa_s0_c63_n334_s;
                stage1_col63[15] = fa_s0_c63_n335_s;
                stage1_col63[16] = fa_s0_c63_n336_s;
                stage1_col63[17] = fa_s0_c63_n337_s;
                stage1_col63[18] = fa_s0_c63_n338_s;
                stage1_col63[19] = fa_s0_c63_n339_s;
                stage1_col63[20] = fa_s0_c63_n340_s;
                stage1_col63[21] = stage0_col63[30];
                stage1_col63[22] = stage0_col63[31];
                stage1_col64[0] = fa_s0_c63_n331_c;
                stage1_col64[1] = fa_s0_c63_n332_c;
                stage1_col64[2] = fa_s0_c63_n333_c;
                stage1_col64[3] = fa_s0_c63_n334_c;
                stage1_col64[4] = fa_s0_c63_n335_c;
                stage1_col64[5] = fa_s0_c63_n336_c;
                stage1_col64[6] = fa_s0_c63_n337_c;
                stage1_col64[7] = fa_s0_c63_n338_c;
                stage1_col64[8] = fa_s0_c63_n339_c;
                stage1_col64[9] = fa_s0_c63_n340_c;
                stage1_col64[10] = fa_s0_c64_n341_s;
                stage1_col64[11] = fa_s0_c64_n342_s;
                stage1_col64[12] = fa_s0_c64_n343_s;
                stage1_col64[13] = fa_s0_c64_n344_s;
                stage1_col64[14] = fa_s0_c64_n345_s;
                stage1_col64[15] = fa_s0_c64_n346_s;
                stage1_col64[16] = fa_s0_c64_n347_s;
                stage1_col64[17] = fa_s0_c64_n348_s;
                stage1_col64[18] = fa_s0_c64_n349_s;
                stage1_col64[19] = fa_s0_c64_n350_s;
                stage1_col64[20] = fa_s0_c64_n351_s;
                stage1_col65[0] = fa_s0_c64_n341_c;
                stage1_col65[1] = fa_s0_c64_n342_c;
                stage1_col65[2] = fa_s0_c64_n343_c;
                stage1_col65[3] = fa_s0_c64_n344_c;
                stage1_col65[4] = fa_s0_c64_n345_c;
                stage1_col65[5] = fa_s0_c64_n346_c;
                stage1_col65[6] = fa_s0_c64_n347_c;
                stage1_col65[7] = fa_s0_c64_n348_c;
                stage1_col65[8] = fa_s0_c64_n349_c;
                stage1_col65[9] = fa_s0_c64_n350_c;
                stage1_col65[10] = fa_s0_c64_n351_c;
                stage1_col65[11] = fa_s0_c65_n352_s;
                stage1_col65[12] = fa_s0_c65_n353_s;
                stage1_col65[13] = fa_s0_c65_n354_s;
                stage1_col65[14] = fa_s0_c65_n355_s;
                stage1_col65[15] = fa_s0_c65_n356_s;
                stage1_col65[16] = fa_s0_c65_n357_s;
                stage1_col65[17] = fa_s0_c65_n358_s;
                stage1_col65[18] = fa_s0_c65_n359_s;
                stage1_col65[19] = fa_s0_c65_n360_s;
                stage1_col65[20] = fa_s0_c65_n361_s;
                stage1_col65[21] = stage0_col65[30];
                stage1_col65[22] = stage0_col65[31];
                stage1_col66[0] = fa_s0_c65_n352_c;
                stage1_col66[1] = fa_s0_c65_n353_c;
                stage1_col66[2] = fa_s0_c65_n354_c;
                stage1_col66[3] = fa_s0_c65_n355_c;
                stage1_col66[4] = fa_s0_c65_n356_c;
                stage1_col66[5] = fa_s0_c65_n357_c;
                stage1_col66[6] = fa_s0_c65_n358_c;
                stage1_col66[7] = fa_s0_c65_n359_c;
                stage1_col66[8] = fa_s0_c65_n360_c;
                stage1_col66[9] = fa_s0_c65_n361_c;
                stage1_col66[10] = fa_s0_c66_n362_s;
                stage1_col66[11] = fa_s0_c66_n363_s;
                stage1_col66[12] = fa_s0_c66_n364_s;
                stage1_col66[13] = fa_s0_c66_n365_s;
                stage1_col66[14] = fa_s0_c66_n366_s;
                stage1_col66[15] = fa_s0_c66_n367_s;
                stage1_col66[16] = fa_s0_c66_n368_s;
                stage1_col66[17] = fa_s0_c66_n369_s;
                stage1_col66[18] = fa_s0_c66_n370_s;
                stage1_col66[19] = fa_s0_c66_n371_s;
                stage1_col66[20] = fa_s0_c66_n372_s;
                stage1_col67[0] = fa_s0_c66_n362_c;
                stage1_col67[1] = fa_s0_c66_n363_c;
                stage1_col67[2] = fa_s0_c66_n364_c;
                stage1_col67[3] = fa_s0_c66_n365_c;
                stage1_col67[4] = fa_s0_c66_n366_c;
                stage1_col67[5] = fa_s0_c66_n367_c;
                stage1_col67[6] = fa_s0_c66_n368_c;
                stage1_col67[7] = fa_s0_c66_n369_c;
                stage1_col67[8] = fa_s0_c66_n370_c;
                stage1_col67[9] = fa_s0_c66_n371_c;
                stage1_col67[10] = fa_s0_c66_n372_c;
                stage1_col67[11] = fa_s0_c67_n373_s;
                stage1_col67[12] = fa_s0_c67_n374_s;
                stage1_col67[13] = fa_s0_c67_n375_s;
                stage1_col67[14] = fa_s0_c67_n376_s;
                stage1_col67[15] = fa_s0_c67_n377_s;
                stage1_col67[16] = fa_s0_c67_n378_s;
                stage1_col67[17] = fa_s0_c67_n379_s;
                stage1_col67[18] = fa_s0_c67_n380_s;
                stage1_col67[19] = fa_s0_c67_n381_s;
                stage1_col67[20] = fa_s0_c67_n382_s;
                stage1_col67[21] = stage0_col67[30];
                stage1_col67[22] = stage0_col67[31];
                stage1_col68[0] = fa_s0_c67_n373_c;
                stage1_col68[1] = fa_s0_c67_n374_c;
                stage1_col68[2] = fa_s0_c67_n375_c;
                stage1_col68[3] = fa_s0_c67_n376_c;
                stage1_col68[4] = fa_s0_c67_n377_c;
                stage1_col68[5] = fa_s0_c67_n378_c;
                stage1_col68[6] = fa_s0_c67_n379_c;
                stage1_col68[7] = fa_s0_c67_n380_c;
                stage1_col68[8] = fa_s0_c67_n381_c;
                stage1_col68[9] = fa_s0_c67_n382_c;
                stage1_col68[10] = fa_s0_c68_n383_s;
                stage1_col68[11] = fa_s0_c68_n384_s;
                stage1_col68[12] = fa_s0_c68_n385_s;
                stage1_col68[13] = fa_s0_c68_n386_s;
                stage1_col68[14] = fa_s0_c68_n387_s;
                stage1_col68[15] = fa_s0_c68_n388_s;
                stage1_col68[16] = fa_s0_c68_n389_s;
                stage1_col68[17] = fa_s0_c68_n390_s;
                stage1_col68[18] = fa_s0_c68_n391_s;
                stage1_col68[19] = fa_s0_c68_n392_s;
                stage1_col68[20] = fa_s0_c68_n393_s;
                stage1_col69[0] = fa_s0_c68_n383_c;
                stage1_col69[1] = fa_s0_c68_n384_c;
                stage1_col69[2] = fa_s0_c68_n385_c;
                stage1_col69[3] = fa_s0_c68_n386_c;
                stage1_col69[4] = fa_s0_c68_n387_c;
                stage1_col69[5] = fa_s0_c68_n388_c;
                stage1_col69[6] = fa_s0_c68_n389_c;
                stage1_col69[7] = fa_s0_c68_n390_c;
                stage1_col69[8] = fa_s0_c68_n391_c;
                stage1_col69[9] = fa_s0_c68_n392_c;
                stage1_col69[10] = fa_s0_c68_n393_c;
                stage1_col69[11] = fa_s0_c69_n394_s;
                stage1_col69[12] = fa_s0_c69_n395_s;
                stage1_col69[13] = fa_s0_c69_n396_s;
                stage1_col69[14] = fa_s0_c69_n397_s;
                stage1_col69[15] = fa_s0_c69_n398_s;
                stage1_col69[16] = fa_s0_c69_n399_s;
                stage1_col69[17] = fa_s0_c69_n400_s;
                stage1_col69[18] = fa_s0_c69_n401_s;
                stage1_col69[19] = fa_s0_c69_n402_s;
                stage1_col69[20] = fa_s0_c69_n403_s;
                stage1_col69[21] = stage0_col69[30];
                stage1_col69[22] = stage0_col69[31];
                stage1_col70[0] = fa_s0_c69_n394_c;
                stage1_col70[1] = fa_s0_c69_n395_c;
                stage1_col70[2] = fa_s0_c69_n396_c;
                stage1_col70[3] = fa_s0_c69_n397_c;
                stage1_col70[4] = fa_s0_c69_n398_c;
                stage1_col70[5] = fa_s0_c69_n399_c;
                stage1_col70[6] = fa_s0_c69_n400_c;
                stage1_col70[7] = fa_s0_c69_n401_c;
                stage1_col70[8] = fa_s0_c69_n402_c;
                stage1_col70[9] = fa_s0_c69_n403_c;
                stage1_col70[10] = fa_s0_c70_n404_s;
                stage1_col70[11] = fa_s0_c70_n405_s;
                stage1_col70[12] = fa_s0_c70_n406_s;
                stage1_col70[13] = fa_s0_c70_n407_s;
                stage1_col70[14] = fa_s0_c70_n408_s;
                stage1_col70[15] = fa_s0_c70_n409_s;
                stage1_col70[16] = fa_s0_c70_n410_s;
                stage1_col70[17] = fa_s0_c70_n411_s;
                stage1_col70[18] = fa_s0_c70_n412_s;
                stage1_col70[19] = fa_s0_c70_n413_s;
                stage1_col70[20] = fa_s0_c70_n414_s;
                stage1_col71[0] = fa_s0_c70_n404_c;
                stage1_col71[1] = fa_s0_c70_n405_c;
                stage1_col71[2] = fa_s0_c70_n406_c;
                stage1_col71[3] = fa_s0_c70_n407_c;
                stage1_col71[4] = fa_s0_c70_n408_c;
                stage1_col71[5] = fa_s0_c70_n409_c;
                stage1_col71[6] = fa_s0_c70_n410_c;
                stage1_col71[7] = fa_s0_c70_n411_c;
                stage1_col71[8] = fa_s0_c70_n412_c;
                stage1_col71[9] = fa_s0_c70_n413_c;
                stage1_col71[10] = fa_s0_c70_n414_c;
                stage1_col71[11] = fa_s0_c71_n415_s;
                stage1_col71[12] = fa_s0_c71_n416_s;
                stage1_col71[13] = fa_s0_c71_n417_s;
                stage1_col71[14] = fa_s0_c71_n418_s;
                stage1_col71[15] = fa_s0_c71_n419_s;
                stage1_col71[16] = fa_s0_c71_n420_s;
                stage1_col71[17] = fa_s0_c71_n421_s;
                stage1_col71[18] = fa_s0_c71_n422_s;
                stage1_col71[19] = fa_s0_c71_n423_s;
                stage1_col71[20] = fa_s0_c71_n424_s;
                stage1_col71[21] = stage0_col71[30];
                stage1_col71[22] = stage0_col71[31];
                stage1_col72[0] = fa_s0_c71_n415_c;
                stage1_col72[1] = fa_s0_c71_n416_c;
                stage1_col72[2] = fa_s0_c71_n417_c;
                stage1_col72[3] = fa_s0_c71_n418_c;
                stage1_col72[4] = fa_s0_c71_n419_c;
                stage1_col72[5] = fa_s0_c71_n420_c;
                stage1_col72[6] = fa_s0_c71_n421_c;
                stage1_col72[7] = fa_s0_c71_n422_c;
                stage1_col72[8] = fa_s0_c71_n423_c;
                stage1_col72[9] = fa_s0_c71_n424_c;
                stage1_col72[10] = fa_s0_c72_n425_s;
                stage1_col72[11] = fa_s0_c72_n426_s;
                stage1_col72[12] = fa_s0_c72_n427_s;
                stage1_col72[13] = fa_s0_c72_n428_s;
                stage1_col72[14] = fa_s0_c72_n429_s;
                stage1_col72[15] = fa_s0_c72_n430_s;
                stage1_col72[16] = fa_s0_c72_n431_s;
                stage1_col72[17] = fa_s0_c72_n432_s;
                stage1_col72[18] = fa_s0_c72_n433_s;
                stage1_col72[19] = fa_s0_c72_n434_s;
                stage1_col72[20] = fa_s0_c72_n435_s;
                stage1_col73[0] = fa_s0_c72_n425_c;
                stage1_col73[1] = fa_s0_c72_n426_c;
                stage1_col73[2] = fa_s0_c72_n427_c;
                stage1_col73[3] = fa_s0_c72_n428_c;
                stage1_col73[4] = fa_s0_c72_n429_c;
                stage1_col73[5] = fa_s0_c72_n430_c;
                stage1_col73[6] = fa_s0_c72_n431_c;
                stage1_col73[7] = fa_s0_c72_n432_c;
                stage1_col73[8] = fa_s0_c72_n433_c;
                stage1_col73[9] = fa_s0_c72_n434_c;
                stage1_col73[10] = fa_s0_c72_n435_c;
                stage1_col73[11] = fa_s0_c73_n436_s;
                stage1_col73[12] = fa_s0_c73_n437_s;
                stage1_col73[13] = fa_s0_c73_n438_s;
                stage1_col73[14] = fa_s0_c73_n439_s;
                stage1_col73[15] = fa_s0_c73_n440_s;
                stage1_col73[16] = fa_s0_c73_n441_s;
                stage1_col73[17] = fa_s0_c73_n442_s;
                stage1_col73[18] = fa_s0_c73_n443_s;
                stage1_col73[19] = fa_s0_c73_n444_s;
                stage1_col73[20] = fa_s0_c73_n445_s;
                stage1_col73[21] = stage0_col73[30];
                stage1_col73[22] = stage0_col73[31];
                stage1_col74[0] = fa_s0_c73_n436_c;
                stage1_col74[1] = fa_s0_c73_n437_c;
                stage1_col74[2] = fa_s0_c73_n438_c;
                stage1_col74[3] = fa_s0_c73_n439_c;
                stage1_col74[4] = fa_s0_c73_n440_c;
                stage1_col74[5] = fa_s0_c73_n441_c;
                stage1_col74[6] = fa_s0_c73_n442_c;
                stage1_col74[7] = fa_s0_c73_n443_c;
                stage1_col74[8] = fa_s0_c73_n444_c;
                stage1_col74[9] = fa_s0_c73_n445_c;
                stage1_col74[10] = fa_s0_c74_n446_s;
                stage1_col74[11] = fa_s0_c74_n447_s;
                stage1_col74[12] = fa_s0_c74_n448_s;
                stage1_col74[13] = fa_s0_c74_n449_s;
                stage1_col74[14] = fa_s0_c74_n450_s;
                stage1_col74[15] = fa_s0_c74_n451_s;
                stage1_col74[16] = fa_s0_c74_n452_s;
                stage1_col74[17] = fa_s0_c74_n453_s;
                stage1_col74[18] = fa_s0_c74_n454_s;
                stage1_col74[19] = fa_s0_c74_n455_s;
                stage1_col74[20] = fa_s0_c74_n456_s;
                stage1_col75[0] = fa_s0_c74_n446_c;
                stage1_col75[1] = fa_s0_c74_n447_c;
                stage1_col75[2] = fa_s0_c74_n448_c;
                stage1_col75[3] = fa_s0_c74_n449_c;
                stage1_col75[4] = fa_s0_c74_n450_c;
                stage1_col75[5] = fa_s0_c74_n451_c;
                stage1_col75[6] = fa_s0_c74_n452_c;
                stage1_col75[7] = fa_s0_c74_n453_c;
                stage1_col75[8] = fa_s0_c74_n454_c;
                stage1_col75[9] = fa_s0_c74_n455_c;
                stage1_col75[10] = fa_s0_c74_n456_c;
                stage1_col75[11] = fa_s0_c75_n457_s;
                stage1_col75[12] = fa_s0_c75_n458_s;
                stage1_col75[13] = fa_s0_c75_n459_s;
                stage1_col75[14] = fa_s0_c75_n460_s;
                stage1_col75[15] = fa_s0_c75_n461_s;
                stage1_col75[16] = fa_s0_c75_n462_s;
                stage1_col75[17] = fa_s0_c75_n463_s;
                stage1_col75[18] = fa_s0_c75_n464_s;
                stage1_col75[19] = fa_s0_c75_n465_s;
                stage1_col75[20] = fa_s0_c75_n466_s;
                stage1_col75[21] = stage0_col75[30];
                stage1_col75[22] = stage0_col75[31];
                stage1_col76[0] = fa_s0_c75_n457_c;
                stage1_col76[1] = fa_s0_c75_n458_c;
                stage1_col76[2] = fa_s0_c75_n459_c;
                stage1_col76[3] = fa_s0_c75_n460_c;
                stage1_col76[4] = fa_s0_c75_n461_c;
                stage1_col76[5] = fa_s0_c75_n462_c;
                stage1_col76[6] = fa_s0_c75_n463_c;
                stage1_col76[7] = fa_s0_c75_n464_c;
                stage1_col76[8] = fa_s0_c75_n465_c;
                stage1_col76[9] = fa_s0_c75_n466_c;
                stage1_col76[10] = fa_s0_c76_n467_s;
                stage1_col76[11] = fa_s0_c76_n468_s;
                stage1_col76[12] = fa_s0_c76_n469_s;
                stage1_col76[13] = fa_s0_c76_n470_s;
                stage1_col76[14] = fa_s0_c76_n471_s;
                stage1_col76[15] = fa_s0_c76_n472_s;
                stage1_col76[16] = fa_s0_c76_n473_s;
                stage1_col76[17] = fa_s0_c76_n474_s;
                stage1_col76[18] = fa_s0_c76_n475_s;
                stage1_col76[19] = fa_s0_c76_n476_s;
                stage1_col76[20] = fa_s0_c76_n477_s;
                stage1_col77[0] = fa_s0_c76_n467_c;
                stage1_col77[1] = fa_s0_c76_n468_c;
                stage1_col77[2] = fa_s0_c76_n469_c;
                stage1_col77[3] = fa_s0_c76_n470_c;
                stage1_col77[4] = fa_s0_c76_n471_c;
                stage1_col77[5] = fa_s0_c76_n472_c;
                stage1_col77[6] = fa_s0_c76_n473_c;
                stage1_col77[7] = fa_s0_c76_n474_c;
                stage1_col77[8] = fa_s0_c76_n475_c;
                stage1_col77[9] = fa_s0_c76_n476_c;
                stage1_col77[10] = fa_s0_c76_n477_c;
                stage1_col77[11] = fa_s0_c77_n478_s;
                stage1_col77[12] = fa_s0_c77_n479_s;
                stage1_col77[13] = fa_s0_c77_n480_s;
                stage1_col77[14] = fa_s0_c77_n481_s;
                stage1_col77[15] = fa_s0_c77_n482_s;
                stage1_col77[16] = fa_s0_c77_n483_s;
                stage1_col77[17] = fa_s0_c77_n484_s;
                stage1_col77[18] = fa_s0_c77_n485_s;
                stage1_col77[19] = fa_s0_c77_n486_s;
                stage1_col77[20] = fa_s0_c77_n487_s;
                stage1_col77[21] = stage0_col77[30];
                stage1_col77[22] = stage0_col77[31];
                stage1_col78[0] = fa_s0_c77_n478_c;
                stage1_col78[1] = fa_s0_c77_n479_c;
                stage1_col78[2] = fa_s0_c77_n480_c;
                stage1_col78[3] = fa_s0_c77_n481_c;
                stage1_col78[4] = fa_s0_c77_n482_c;
                stage1_col78[5] = fa_s0_c77_n483_c;
                stage1_col78[6] = fa_s0_c77_n484_c;
                stage1_col78[7] = fa_s0_c77_n485_c;
                stage1_col78[8] = fa_s0_c77_n486_c;
                stage1_col78[9] = fa_s0_c77_n487_c;
                stage1_col78[10] = fa_s0_c78_n488_s;
                stage1_col78[11] = fa_s0_c78_n489_s;
                stage1_col78[12] = fa_s0_c78_n490_s;
                stage1_col78[13] = fa_s0_c78_n491_s;
                stage1_col78[14] = fa_s0_c78_n492_s;
                stage1_col78[15] = fa_s0_c78_n493_s;
                stage1_col78[16] = fa_s0_c78_n494_s;
                stage1_col78[17] = fa_s0_c78_n495_s;
                stage1_col78[18] = fa_s0_c78_n496_s;
                stage1_col78[19] = fa_s0_c78_n497_s;
                stage1_col78[20] = fa_s0_c78_n498_s;
                stage1_col79[0] = fa_s0_c78_n488_c;
                stage1_col79[1] = fa_s0_c78_n489_c;
                stage1_col79[2] = fa_s0_c78_n490_c;
                stage1_col79[3] = fa_s0_c78_n491_c;
                stage1_col79[4] = fa_s0_c78_n492_c;
                stage1_col79[5] = fa_s0_c78_n493_c;
                stage1_col79[6] = fa_s0_c78_n494_c;
                stage1_col79[7] = fa_s0_c78_n495_c;
                stage1_col79[8] = fa_s0_c78_n496_c;
                stage1_col79[9] = fa_s0_c78_n497_c;
                stage1_col79[10] = fa_s0_c78_n498_c;
                stage1_col79[11] = fa_s0_c79_n499_s;
                stage1_col79[12] = fa_s0_c79_n500_s;
                stage1_col79[13] = fa_s0_c79_n501_s;
                stage1_col79[14] = fa_s0_c79_n502_s;
                stage1_col79[15] = fa_s0_c79_n503_s;
                stage1_col79[16] = fa_s0_c79_n504_s;
                stage1_col79[17] = fa_s0_c79_n505_s;
                stage1_col79[18] = fa_s0_c79_n506_s;
                stage1_col79[19] = fa_s0_c79_n507_s;
                stage1_col79[20] = fa_s0_c79_n508_s;
                stage1_col79[21] = stage0_col79[30];
                stage1_col79[22] = stage0_col79[31];
                stage1_col80[0] = fa_s0_c79_n499_c;
                stage1_col80[1] = fa_s0_c79_n500_c;
                stage1_col80[2] = fa_s0_c79_n501_c;
                stage1_col80[3] = fa_s0_c79_n502_c;
                stage1_col80[4] = fa_s0_c79_n503_c;
                stage1_col80[5] = fa_s0_c79_n504_c;
                stage1_col80[6] = fa_s0_c79_n505_c;
                stage1_col80[7] = fa_s0_c79_n506_c;
                stage1_col80[8] = fa_s0_c79_n507_c;
                stage1_col80[9] = fa_s0_c79_n508_c;
                stage1_col80[10] = fa_s0_c80_n509_s;
                stage1_col80[11] = fa_s0_c80_n510_s;
                stage1_col80[12] = fa_s0_c80_n511_s;
                stage1_col80[13] = fa_s0_c80_n512_s;
                stage1_col80[14] = fa_s0_c80_n513_s;
                stage1_col80[15] = fa_s0_c80_n514_s;
                stage1_col80[16] = fa_s0_c80_n515_s;
                stage1_col80[17] = fa_s0_c80_n516_s;
                stage1_col80[18] = fa_s0_c80_n517_s;
                stage1_col80[19] = fa_s0_c80_n518_s;
                stage1_col80[20] = fa_s0_c80_n519_s;
                stage1_col81[0] = fa_s0_c80_n509_c;
                stage1_col81[1] = fa_s0_c80_n510_c;
                stage1_col81[2] = fa_s0_c80_n511_c;
                stage1_col81[3] = fa_s0_c80_n512_c;
                stage1_col81[4] = fa_s0_c80_n513_c;
                stage1_col81[5] = fa_s0_c80_n514_c;
                stage1_col81[6] = fa_s0_c80_n515_c;
                stage1_col81[7] = fa_s0_c80_n516_c;
                stage1_col81[8] = fa_s0_c80_n517_c;
                stage1_col81[9] = fa_s0_c80_n518_c;
                stage1_col81[10] = fa_s0_c80_n519_c;
                stage1_col81[11] = fa_s0_c81_n520_s;
                stage1_col81[12] = fa_s0_c81_n521_s;
                stage1_col81[13] = fa_s0_c81_n522_s;
                stage1_col81[14] = fa_s0_c81_n523_s;
                stage1_col81[15] = fa_s0_c81_n524_s;
                stage1_col81[16] = fa_s0_c81_n525_s;
                stage1_col81[17] = fa_s0_c81_n526_s;
                stage1_col81[18] = fa_s0_c81_n527_s;
                stage1_col81[19] = fa_s0_c81_n528_s;
                stage1_col81[20] = fa_s0_c81_n529_s;
                stage1_col81[21] = stage0_col81[30];
                stage1_col81[22] = stage0_col81[31];
                stage1_col82[0] = fa_s0_c81_n520_c;
                stage1_col82[1] = fa_s0_c81_n521_c;
                stage1_col82[2] = fa_s0_c81_n522_c;
                stage1_col82[3] = fa_s0_c81_n523_c;
                stage1_col82[4] = fa_s0_c81_n524_c;
                stage1_col82[5] = fa_s0_c81_n525_c;
                stage1_col82[6] = fa_s0_c81_n526_c;
                stage1_col82[7] = fa_s0_c81_n527_c;
                stage1_col82[8] = fa_s0_c81_n528_c;
                stage1_col82[9] = fa_s0_c81_n529_c;
                stage1_col82[10] = fa_s0_c82_n530_s;
                stage1_col82[11] = fa_s0_c82_n531_s;
                stage1_col82[12] = fa_s0_c82_n532_s;
                stage1_col82[13] = fa_s0_c82_n533_s;
                stage1_col82[14] = fa_s0_c82_n534_s;
                stage1_col82[15] = fa_s0_c82_n535_s;
                stage1_col82[16] = fa_s0_c82_n536_s;
                stage1_col82[17] = fa_s0_c82_n537_s;
                stage1_col82[18] = fa_s0_c82_n538_s;
                stage1_col82[19] = fa_s0_c82_n539_s;
                stage1_col82[20] = fa_s0_c82_n540_s;
                stage1_col83[0] = fa_s0_c82_n530_c;
                stage1_col83[1] = fa_s0_c82_n531_c;
                stage1_col83[2] = fa_s0_c82_n532_c;
                stage1_col83[3] = fa_s0_c82_n533_c;
                stage1_col83[4] = fa_s0_c82_n534_c;
                stage1_col83[5] = fa_s0_c82_n535_c;
                stage1_col83[6] = fa_s0_c82_n536_c;
                stage1_col83[7] = fa_s0_c82_n537_c;
                stage1_col83[8] = fa_s0_c82_n538_c;
                stage1_col83[9] = fa_s0_c82_n539_c;
                stage1_col83[10] = fa_s0_c82_n540_c;
                stage1_col83[11] = fa_s0_c83_n541_s;
                stage1_col83[12] = fa_s0_c83_n542_s;
                stage1_col83[13] = fa_s0_c83_n543_s;
                stage1_col83[14] = fa_s0_c83_n544_s;
                stage1_col83[15] = fa_s0_c83_n545_s;
                stage1_col83[16] = fa_s0_c83_n546_s;
                stage1_col83[17] = fa_s0_c83_n547_s;
                stage1_col83[18] = fa_s0_c83_n548_s;
                stage1_col83[19] = fa_s0_c83_n549_s;
                stage1_col83[20] = fa_s0_c83_n550_s;
                stage1_col83[21] = stage0_col83[30];
                stage1_col83[22] = stage0_col83[31];
                stage1_col84[0] = fa_s0_c83_n541_c;
                stage1_col84[1] = fa_s0_c83_n542_c;
                stage1_col84[2] = fa_s0_c83_n543_c;
                stage1_col84[3] = fa_s0_c83_n544_c;
                stage1_col84[4] = fa_s0_c83_n545_c;
                stage1_col84[5] = fa_s0_c83_n546_c;
                stage1_col84[6] = fa_s0_c83_n547_c;
                stage1_col84[7] = fa_s0_c83_n548_c;
                stage1_col84[8] = fa_s0_c83_n549_c;
                stage1_col84[9] = fa_s0_c83_n550_c;
                stage1_col84[10] = fa_s0_c84_n551_s;
                stage1_col84[11] = fa_s0_c84_n552_s;
                stage1_col84[12] = fa_s0_c84_n553_s;
                stage1_col84[13] = fa_s0_c84_n554_s;
                stage1_col84[14] = fa_s0_c84_n555_s;
                stage1_col84[15] = fa_s0_c84_n556_s;
                stage1_col84[16] = fa_s0_c84_n557_s;
                stage1_col84[17] = fa_s0_c84_n558_s;
                stage1_col84[18] = fa_s0_c84_n559_s;
                stage1_col84[19] = fa_s0_c84_n560_s;
                stage1_col84[20] = fa_s0_c84_n561_s;
                stage1_col85[0] = fa_s0_c84_n551_c;
                stage1_col85[1] = fa_s0_c84_n552_c;
                stage1_col85[2] = fa_s0_c84_n553_c;
                stage1_col85[3] = fa_s0_c84_n554_c;
                stage1_col85[4] = fa_s0_c84_n555_c;
                stage1_col85[5] = fa_s0_c84_n556_c;
                stage1_col85[6] = fa_s0_c84_n557_c;
                stage1_col85[7] = fa_s0_c84_n558_c;
                stage1_col85[8] = fa_s0_c84_n559_c;
                stage1_col85[9] = fa_s0_c84_n560_c;
                stage1_col85[10] = fa_s0_c84_n561_c;
                stage1_col85[11] = fa_s0_c85_n562_s;
                stage1_col85[12] = fa_s0_c85_n563_s;
                stage1_col85[13] = fa_s0_c85_n564_s;
                stage1_col85[14] = fa_s0_c85_n565_s;
                stage1_col85[15] = fa_s0_c85_n566_s;
                stage1_col85[16] = fa_s0_c85_n567_s;
                stage1_col85[17] = fa_s0_c85_n568_s;
                stage1_col85[18] = fa_s0_c85_n569_s;
                stage1_col85[19] = fa_s0_c85_n570_s;
                stage1_col85[20] = fa_s0_c85_n571_s;
                stage1_col85[21] = stage0_col85[30];
                stage1_col85[22] = stage0_col85[31];
                stage1_col86[0] = fa_s0_c85_n562_c;
                stage1_col86[1] = fa_s0_c85_n563_c;
                stage1_col86[2] = fa_s0_c85_n564_c;
                stage1_col86[3] = fa_s0_c85_n565_c;
                stage1_col86[4] = fa_s0_c85_n566_c;
                stage1_col86[5] = fa_s0_c85_n567_c;
                stage1_col86[6] = fa_s0_c85_n568_c;
                stage1_col86[7] = fa_s0_c85_n569_c;
                stage1_col86[8] = fa_s0_c85_n570_c;
                stage1_col86[9] = fa_s0_c85_n571_c;
                stage1_col86[10] = fa_s0_c86_n572_s;
                stage1_col86[11] = fa_s0_c86_n573_s;
                stage1_col86[12] = fa_s0_c86_n574_s;
                stage1_col86[13] = fa_s0_c86_n575_s;
                stage1_col86[14] = fa_s0_c86_n576_s;
                stage1_col86[15] = fa_s0_c86_n577_s;
                stage1_col86[16] = fa_s0_c86_n578_s;
                stage1_col86[17] = fa_s0_c86_n579_s;
                stage1_col86[18] = fa_s0_c86_n580_s;
                stage1_col86[19] = fa_s0_c86_n581_s;
                stage1_col86[20] = fa_s0_c86_n582_s;
                stage1_col87[0] = fa_s0_c86_n572_c;
                stage1_col87[1] = fa_s0_c86_n573_c;
                stage1_col87[2] = fa_s0_c86_n574_c;
                stage1_col87[3] = fa_s0_c86_n575_c;
                stage1_col87[4] = fa_s0_c86_n576_c;
                stage1_col87[5] = fa_s0_c86_n577_c;
                stage1_col87[6] = fa_s0_c86_n578_c;
                stage1_col87[7] = fa_s0_c86_n579_c;
                stage1_col87[8] = fa_s0_c86_n580_c;
                stage1_col87[9] = fa_s0_c86_n581_c;
                stage1_col87[10] = fa_s0_c86_n582_c;
                stage1_col87[11] = fa_s0_c87_n583_s;
                stage1_col87[12] = fa_s0_c87_n584_s;
                stage1_col87[13] = fa_s0_c87_n585_s;
                stage1_col87[14] = fa_s0_c87_n586_s;
                stage1_col87[15] = fa_s0_c87_n587_s;
                stage1_col87[16] = fa_s0_c87_n588_s;
                stage1_col87[17] = fa_s0_c87_n589_s;
                stage1_col87[18] = fa_s0_c87_n590_s;
                stage1_col87[19] = fa_s0_c87_n591_s;
                stage1_col87[20] = fa_s0_c87_n592_s;
                stage1_col87[21] = stage0_col87[30];
                stage1_col87[22] = stage0_col87[31];
                stage1_col88[0] = fa_s0_c87_n583_c;
                stage1_col88[1] = fa_s0_c87_n584_c;
                stage1_col88[2] = fa_s0_c87_n585_c;
                stage1_col88[3] = fa_s0_c87_n586_c;
                stage1_col88[4] = fa_s0_c87_n587_c;
                stage1_col88[5] = fa_s0_c87_n588_c;
                stage1_col88[6] = fa_s0_c87_n589_c;
                stage1_col88[7] = fa_s0_c87_n590_c;
                stage1_col88[8] = fa_s0_c87_n591_c;
                stage1_col88[9] = fa_s0_c87_n592_c;
                stage1_col88[10] = fa_s0_c88_n593_s;
                stage1_col88[11] = fa_s0_c88_n594_s;
                stage1_col88[12] = fa_s0_c88_n595_s;
                stage1_col88[13] = fa_s0_c88_n596_s;
                stage1_col88[14] = fa_s0_c88_n597_s;
                stage1_col88[15] = fa_s0_c88_n598_s;
                stage1_col88[16] = fa_s0_c88_n599_s;
                stage1_col88[17] = fa_s0_c88_n600_s;
                stage1_col88[18] = fa_s0_c88_n601_s;
                stage1_col88[19] = fa_s0_c88_n602_s;
                stage1_col88[20] = fa_s0_c88_n603_s;
                stage1_col89[0] = fa_s0_c88_n593_c;
                stage1_col89[1] = fa_s0_c88_n594_c;
                stage1_col89[2] = fa_s0_c88_n595_c;
                stage1_col89[3] = fa_s0_c88_n596_c;
                stage1_col89[4] = fa_s0_c88_n597_c;
                stage1_col89[5] = fa_s0_c88_n598_c;
                stage1_col89[6] = fa_s0_c88_n599_c;
                stage1_col89[7] = fa_s0_c88_n600_c;
                stage1_col89[8] = fa_s0_c88_n601_c;
                stage1_col89[9] = fa_s0_c88_n602_c;
                stage1_col89[10] = fa_s0_c88_n603_c;
                stage1_col89[11] = fa_s0_c89_n604_s;
                stage1_col89[12] = fa_s0_c89_n605_s;
                stage1_col89[13] = fa_s0_c89_n606_s;
                stage1_col89[14] = fa_s0_c89_n607_s;
                stage1_col89[15] = fa_s0_c89_n608_s;
                stage1_col89[16] = fa_s0_c89_n609_s;
                stage1_col89[17] = fa_s0_c89_n610_s;
                stage1_col89[18] = fa_s0_c89_n611_s;
                stage1_col89[19] = fa_s0_c89_n612_s;
                stage1_col89[20] = fa_s0_c89_n613_s;
                stage1_col89[21] = stage0_col89[30];
                stage1_col89[22] = stage0_col89[31];
                stage1_col90[0] = fa_s0_c89_n604_c;
                stage1_col90[1] = fa_s0_c89_n605_c;
                stage1_col90[2] = fa_s0_c89_n606_c;
                stage1_col90[3] = fa_s0_c89_n607_c;
                stage1_col90[4] = fa_s0_c89_n608_c;
                stage1_col90[5] = fa_s0_c89_n609_c;
                stage1_col90[6] = fa_s0_c89_n610_c;
                stage1_col90[7] = fa_s0_c89_n611_c;
                stage1_col90[8] = fa_s0_c89_n612_c;
                stage1_col90[9] = fa_s0_c89_n613_c;
                stage1_col90[10] = fa_s0_c90_n614_s;
                stage1_col90[11] = fa_s0_c90_n615_s;
                stage1_col90[12] = fa_s0_c90_n616_s;
                stage1_col90[13] = fa_s0_c90_n617_s;
                stage1_col90[14] = fa_s0_c90_n618_s;
                stage1_col90[15] = fa_s0_c90_n619_s;
                stage1_col90[16] = fa_s0_c90_n620_s;
                stage1_col90[17] = fa_s0_c90_n621_s;
                stage1_col90[18] = fa_s0_c90_n622_s;
                stage1_col90[19] = fa_s0_c90_n623_s;
                stage1_col90[20] = fa_s0_c90_n624_s;
                stage1_col91[0] = fa_s0_c90_n614_c;
                stage1_col91[1] = fa_s0_c90_n615_c;
                stage1_col91[2] = fa_s0_c90_n616_c;
                stage1_col91[3] = fa_s0_c90_n617_c;
                stage1_col91[4] = fa_s0_c90_n618_c;
                stage1_col91[5] = fa_s0_c90_n619_c;
                stage1_col91[6] = fa_s0_c90_n620_c;
                stage1_col91[7] = fa_s0_c90_n621_c;
                stage1_col91[8] = fa_s0_c90_n622_c;
                stage1_col91[9] = fa_s0_c90_n623_c;
                stage1_col91[10] = fa_s0_c90_n624_c;
                stage1_col91[11] = fa_s0_c91_n625_s;
                stage1_col91[12] = fa_s0_c91_n626_s;
                stage1_col91[13] = fa_s0_c91_n627_s;
                stage1_col91[14] = fa_s0_c91_n628_s;
                stage1_col91[15] = fa_s0_c91_n629_s;
                stage1_col91[16] = fa_s0_c91_n630_s;
                stage1_col91[17] = fa_s0_c91_n631_s;
                stage1_col91[18] = fa_s0_c91_n632_s;
                stage1_col91[19] = fa_s0_c91_n633_s;
                stage1_col91[20] = fa_s0_c91_n634_s;
                stage1_col91[21] = stage0_col91[30];
                stage1_col91[22] = stage0_col91[31];
                stage1_col92[0] = fa_s0_c91_n625_c;
                stage1_col92[1] = fa_s0_c91_n626_c;
                stage1_col92[2] = fa_s0_c91_n627_c;
                stage1_col92[3] = fa_s0_c91_n628_c;
                stage1_col92[4] = fa_s0_c91_n629_c;
                stage1_col92[5] = fa_s0_c91_n630_c;
                stage1_col92[6] = fa_s0_c91_n631_c;
                stage1_col92[7] = fa_s0_c91_n632_c;
                stage1_col92[8] = fa_s0_c91_n633_c;
                stage1_col92[9] = fa_s0_c91_n634_c;
                stage1_col92[10] = fa_s0_c92_n635_s;
                stage1_col92[11] = fa_s0_c92_n636_s;
                stage1_col92[12] = fa_s0_c92_n637_s;
                stage1_col92[13] = fa_s0_c92_n638_s;
                stage1_col92[14] = fa_s0_c92_n639_s;
                stage1_col92[15] = fa_s0_c92_n640_s;
                stage1_col92[16] = fa_s0_c92_n641_s;
                stage1_col92[17] = fa_s0_c92_n642_s;
                stage1_col92[18] = fa_s0_c92_n643_s;
                stage1_col92[19] = fa_s0_c92_n644_s;
                stage1_col92[20] = fa_s0_c92_n645_s;
                stage1_col93[0] = fa_s0_c92_n635_c;
                stage1_col93[1] = fa_s0_c92_n636_c;
                stage1_col93[2] = fa_s0_c92_n637_c;
                stage1_col93[3] = fa_s0_c92_n638_c;
                stage1_col93[4] = fa_s0_c92_n639_c;
                stage1_col93[5] = fa_s0_c92_n640_c;
                stage1_col93[6] = fa_s0_c92_n641_c;
                stage1_col93[7] = fa_s0_c92_n642_c;
                stage1_col93[8] = fa_s0_c92_n643_c;
                stage1_col93[9] = fa_s0_c92_n644_c;
                stage1_col93[10] = fa_s0_c92_n645_c;
                stage1_col93[11] = fa_s0_c93_n646_s;
                stage1_col93[12] = fa_s0_c93_n647_s;
                stage1_col93[13] = fa_s0_c93_n648_s;
                stage1_col93[14] = fa_s0_c93_n649_s;
                stage1_col93[15] = fa_s0_c93_n650_s;
                stage1_col93[16] = fa_s0_c93_n651_s;
                stage1_col93[17] = fa_s0_c93_n652_s;
                stage1_col93[18] = fa_s0_c93_n653_s;
                stage1_col93[19] = fa_s0_c93_n654_s;
                stage1_col93[20] = fa_s0_c93_n655_s;
                stage1_col93[21] = stage0_col93[30];
                stage1_col93[22] = stage0_col93[31];
                stage1_col94[0] = fa_s0_c93_n646_c;
                stage1_col94[1] = fa_s0_c93_n647_c;
                stage1_col94[2] = fa_s0_c93_n648_c;
                stage1_col94[3] = fa_s0_c93_n649_c;
                stage1_col94[4] = fa_s0_c93_n650_c;
                stage1_col94[5] = fa_s0_c93_n651_c;
                stage1_col94[6] = fa_s0_c93_n652_c;
                stage1_col94[7] = fa_s0_c93_n653_c;
                stage1_col94[8] = fa_s0_c93_n654_c;
                stage1_col94[9] = fa_s0_c93_n655_c;
                stage1_col94[10] = fa_s0_c94_n656_s;
                stage1_col94[11] = fa_s0_c94_n657_s;
                stage1_col94[12] = fa_s0_c94_n658_s;
                stage1_col94[13] = fa_s0_c94_n659_s;
                stage1_col94[14] = fa_s0_c94_n660_s;
                stage1_col94[15] = fa_s0_c94_n661_s;
                stage1_col94[16] = fa_s0_c94_n662_s;
                stage1_col94[17] = fa_s0_c94_n663_s;
                stage1_col94[18] = fa_s0_c94_n664_s;
                stage1_col94[19] = fa_s0_c94_n665_s;
                stage1_col94[20] = fa_s0_c94_n666_s;
                stage1_col95[0] = fa_s0_c94_n656_c;
                stage1_col95[1] = fa_s0_c94_n657_c;
                stage1_col95[2] = fa_s0_c94_n658_c;
                stage1_col95[3] = fa_s0_c94_n659_c;
                stage1_col95[4] = fa_s0_c94_n660_c;
                stage1_col95[5] = fa_s0_c94_n661_c;
                stage1_col95[6] = fa_s0_c94_n662_c;
                stage1_col95[7] = fa_s0_c94_n663_c;
                stage1_col95[8] = fa_s0_c94_n664_c;
                stage1_col95[9] = fa_s0_c94_n665_c;
                stage1_col95[10] = fa_s0_c94_n666_c;
                stage1_col95[11] = fa_s0_c95_n667_s;
                stage1_col95[12] = fa_s0_c95_n668_s;
                stage1_col95[13] = fa_s0_c95_n669_s;
                stage1_col95[14] = fa_s0_c95_n670_s;
                stage1_col95[15] = fa_s0_c95_n671_s;
                stage1_col95[16] = fa_s0_c95_n672_s;
                stage1_col95[17] = fa_s0_c95_n673_s;
                stage1_col95[18] = fa_s0_c95_n674_s;
                stage1_col95[19] = fa_s0_c95_n675_s;
                stage1_col95[20] = fa_s0_c95_n676_s;
                stage1_col95[21] = stage0_col95[30];
                stage1_col95[22] = stage0_col95[31];
                stage1_col96[0] = fa_s0_c95_n667_c;
                stage1_col96[1] = fa_s0_c95_n668_c;
                stage1_col96[2] = fa_s0_c95_n669_c;
                stage1_col96[3] = fa_s0_c95_n670_c;
                stage1_col96[4] = fa_s0_c95_n671_c;
                stage1_col96[5] = fa_s0_c95_n672_c;
                stage1_col96[6] = fa_s0_c95_n673_c;
                stage1_col96[7] = fa_s0_c95_n674_c;
                stage1_col96[8] = fa_s0_c95_n675_c;
                stage1_col96[9] = fa_s0_c95_n676_c;
                stage1_col96[10] = fa_s0_c96_n677_s;
                stage1_col96[11] = fa_s0_c96_n678_s;
                stage1_col96[12] = fa_s0_c96_n679_s;
                stage1_col96[13] = fa_s0_c96_n680_s;
                stage1_col96[14] = fa_s0_c96_n681_s;
                stage1_col96[15] = fa_s0_c96_n682_s;
                stage1_col96[16] = fa_s0_c96_n683_s;
                stage1_col96[17] = fa_s0_c96_n684_s;
                stage1_col96[18] = fa_s0_c96_n685_s;
                stage1_col96[19] = fa_s0_c96_n686_s;
                stage1_col96[20] = fa_s0_c96_n687_s;
                stage1_col97[0] = fa_s0_c96_n677_c;
                stage1_col97[1] = fa_s0_c96_n678_c;
                stage1_col97[2] = fa_s0_c96_n679_c;
                stage1_col97[3] = fa_s0_c96_n680_c;
                stage1_col97[4] = fa_s0_c96_n681_c;
                stage1_col97[5] = fa_s0_c96_n682_c;
                stage1_col97[6] = fa_s0_c96_n683_c;
                stage1_col97[7] = fa_s0_c96_n684_c;
                stage1_col97[8] = fa_s0_c96_n685_c;
                stage1_col97[9] = fa_s0_c96_n686_c;
                stage1_col97[10] = fa_s0_c96_n687_c;
                stage1_col97[11] = fa_s0_c97_n688_s;
                stage1_col97[12] = fa_s0_c97_n689_s;
                stage1_col97[13] = fa_s0_c97_n690_s;
                stage1_col97[14] = fa_s0_c97_n691_s;
                stage1_col97[15] = fa_s0_c97_n692_s;
                stage1_col97[16] = fa_s0_c97_n693_s;
                stage1_col97[17] = fa_s0_c97_n694_s;
                stage1_col97[18] = fa_s0_c97_n695_s;
                stage1_col97[19] = fa_s0_c97_n696_s;
                stage1_col97[20] = fa_s0_c97_n697_s;
                stage1_col97[21] = stage0_col97[30];
                stage1_col97[22] = stage0_col97[31];
                stage1_col98[0] = fa_s0_c97_n688_c;
                stage1_col98[1] = fa_s0_c97_n689_c;
                stage1_col98[2] = fa_s0_c97_n690_c;
                stage1_col98[3] = fa_s0_c97_n691_c;
                stage1_col98[4] = fa_s0_c97_n692_c;
                stage1_col98[5] = fa_s0_c97_n693_c;
                stage1_col98[6] = fa_s0_c97_n694_c;
                stage1_col98[7] = fa_s0_c97_n695_c;
                stage1_col98[8] = fa_s0_c97_n696_c;
                stage1_col98[9] = fa_s0_c97_n697_c;
                stage1_col98[10] = fa_s0_c98_n698_s;
                stage1_col98[11] = fa_s0_c98_n699_s;
                stage1_col98[12] = fa_s0_c98_n700_s;
                stage1_col98[13] = fa_s0_c98_n701_s;
                stage1_col98[14] = fa_s0_c98_n702_s;
                stage1_col98[15] = fa_s0_c98_n703_s;
                stage1_col98[16] = fa_s0_c98_n704_s;
                stage1_col98[17] = fa_s0_c98_n705_s;
                stage1_col98[18] = fa_s0_c98_n706_s;
                stage1_col98[19] = fa_s0_c98_n707_s;
                stage1_col98[20] = fa_s0_c98_n708_s;
                stage1_col99[0] = fa_s0_c98_n698_c;
                stage1_col99[1] = fa_s0_c98_n699_c;
                stage1_col99[2] = fa_s0_c98_n700_c;
                stage1_col99[3] = fa_s0_c98_n701_c;
                stage1_col99[4] = fa_s0_c98_n702_c;
                stage1_col99[5] = fa_s0_c98_n703_c;
                stage1_col99[6] = fa_s0_c98_n704_c;
                stage1_col99[7] = fa_s0_c98_n705_c;
                stage1_col99[8] = fa_s0_c98_n706_c;
                stage1_col99[9] = fa_s0_c98_n707_c;
                stage1_col99[10] = fa_s0_c98_n708_c;
                stage1_col99[11] = fa_s0_c99_n709_s;
                stage1_col99[12] = fa_s0_c99_n710_s;
                stage1_col99[13] = fa_s0_c99_n711_s;
                stage1_col99[14] = fa_s0_c99_n712_s;
                stage1_col99[15] = fa_s0_c99_n713_s;
                stage1_col99[16] = fa_s0_c99_n714_s;
                stage1_col99[17] = fa_s0_c99_n715_s;
                stage1_col99[18] = fa_s0_c99_n716_s;
                stage1_col99[19] = fa_s0_c99_n717_s;
                stage1_col99[20] = fa_s0_c99_n718_s;
                stage1_col99[21] = stage0_col99[30];
                stage1_col99[22] = stage0_col99[31];
                stage1_col100[0] = fa_s0_c99_n709_c;
                stage1_col100[1] = fa_s0_c99_n710_c;
                stage1_col100[2] = fa_s0_c99_n711_c;
                stage1_col100[3] = fa_s0_c99_n712_c;
                stage1_col100[4] = fa_s0_c99_n713_c;
                stage1_col100[5] = fa_s0_c99_n714_c;
                stage1_col100[6] = fa_s0_c99_n715_c;
                stage1_col100[7] = fa_s0_c99_n716_c;
                stage1_col100[8] = fa_s0_c99_n717_c;
                stage1_col100[9] = fa_s0_c99_n718_c;
                stage1_col100[10] = fa_s0_c100_n719_s;
                stage1_col100[11] = fa_s0_c100_n720_s;
                stage1_col100[12] = fa_s0_c100_n721_s;
                stage1_col100[13] = fa_s0_c100_n722_s;
                stage1_col100[14] = fa_s0_c100_n723_s;
                stage1_col100[15] = fa_s0_c100_n724_s;
                stage1_col100[16] = fa_s0_c100_n725_s;
                stage1_col100[17] = fa_s0_c100_n726_s;
                stage1_col100[18] = fa_s0_c100_n727_s;
                stage1_col100[19] = fa_s0_c100_n728_s;
                stage1_col100[20] = fa_s0_c100_n729_s;
                stage1_col101[0] = fa_s0_c100_n719_c;
                stage1_col101[1] = fa_s0_c100_n720_c;
                stage1_col101[2] = fa_s0_c100_n721_c;
                stage1_col101[3] = fa_s0_c100_n722_c;
                stage1_col101[4] = fa_s0_c100_n723_c;
                stage1_col101[5] = fa_s0_c100_n724_c;
                stage1_col101[6] = fa_s0_c100_n725_c;
                stage1_col101[7] = fa_s0_c100_n726_c;
                stage1_col101[8] = fa_s0_c100_n727_c;
                stage1_col101[9] = fa_s0_c100_n728_c;
                stage1_col101[10] = fa_s0_c100_n729_c;
                stage1_col101[11] = fa_s0_c101_n730_s;
                stage1_col101[12] = fa_s0_c101_n731_s;
                stage1_col101[13] = fa_s0_c101_n732_s;
                stage1_col101[14] = fa_s0_c101_n733_s;
                stage1_col101[15] = fa_s0_c101_n734_s;
                stage1_col101[16] = fa_s0_c101_n735_s;
                stage1_col101[17] = fa_s0_c101_n736_s;
                stage1_col101[18] = fa_s0_c101_n737_s;
                stage1_col101[19] = fa_s0_c101_n738_s;
                stage1_col101[20] = fa_s0_c101_n739_s;
                stage1_col101[21] = stage0_col101[30];
                stage1_col101[22] = stage0_col101[31];
                stage1_col102[0] = fa_s0_c101_n730_c;
                stage1_col102[1] = fa_s0_c101_n731_c;
                stage1_col102[2] = fa_s0_c101_n732_c;
                stage1_col102[3] = fa_s0_c101_n733_c;
                stage1_col102[4] = fa_s0_c101_n734_c;
                stage1_col102[5] = fa_s0_c101_n735_c;
                stage1_col102[6] = fa_s0_c101_n736_c;
                stage1_col102[7] = fa_s0_c101_n737_c;
                stage1_col102[8] = fa_s0_c101_n738_c;
                stage1_col102[9] = fa_s0_c101_n739_c;
                stage1_col102[10] = fa_s0_c102_n740_s;
                stage1_col102[11] = fa_s0_c102_n741_s;
                stage1_col102[12] = fa_s0_c102_n742_s;
                stage1_col102[13] = fa_s0_c102_n743_s;
                stage1_col102[14] = fa_s0_c102_n744_s;
                stage1_col102[15] = fa_s0_c102_n745_s;
                stage1_col102[16] = fa_s0_c102_n746_s;
                stage1_col102[17] = fa_s0_c102_n747_s;
                stage1_col102[18] = fa_s0_c102_n748_s;
                stage1_col102[19] = fa_s0_c102_n749_s;
                stage1_col102[20] = fa_s0_c102_n750_s;
                stage1_col103[0] = fa_s0_c102_n740_c;
                stage1_col103[1] = fa_s0_c102_n741_c;
                stage1_col103[2] = fa_s0_c102_n742_c;
                stage1_col103[3] = fa_s0_c102_n743_c;
                stage1_col103[4] = fa_s0_c102_n744_c;
                stage1_col103[5] = fa_s0_c102_n745_c;
                stage1_col103[6] = fa_s0_c102_n746_c;
                stage1_col103[7] = fa_s0_c102_n747_c;
                stage1_col103[8] = fa_s0_c102_n748_c;
                stage1_col103[9] = fa_s0_c102_n749_c;
                stage1_col103[10] = fa_s0_c102_n750_c;
                stage1_col103[11] = fa_s0_c103_n751_s;
                stage1_col103[12] = fa_s0_c103_n752_s;
                stage1_col103[13] = fa_s0_c103_n753_s;
                stage1_col103[14] = fa_s0_c103_n754_s;
                stage1_col103[15] = fa_s0_c103_n755_s;
                stage1_col103[16] = fa_s0_c103_n756_s;
                stage1_col103[17] = fa_s0_c103_n757_s;
                stage1_col103[18] = fa_s0_c103_n758_s;
                stage1_col103[19] = fa_s0_c103_n759_s;
                stage1_col103[20] = fa_s0_c103_n760_s;
                stage1_col103[21] = stage0_col103[30];
                stage1_col103[22] = stage0_col103[31];
                stage1_col104[0] = fa_s0_c103_n751_c;
                stage1_col104[1] = fa_s0_c103_n752_c;
                stage1_col104[2] = fa_s0_c103_n753_c;
                stage1_col104[3] = fa_s0_c103_n754_c;
                stage1_col104[4] = fa_s0_c103_n755_c;
                stage1_col104[5] = fa_s0_c103_n756_c;
                stage1_col104[6] = fa_s0_c103_n757_c;
                stage1_col104[7] = fa_s0_c103_n758_c;
                stage1_col104[8] = fa_s0_c103_n759_c;
                stage1_col104[9] = fa_s0_c103_n760_c;
                stage1_col104[10] = fa_s0_c104_n761_s;
                stage1_col104[11] = fa_s0_c104_n762_s;
                stage1_col104[12] = fa_s0_c104_n763_s;
                stage1_col104[13] = fa_s0_c104_n764_s;
                stage1_col104[14] = fa_s0_c104_n765_s;
                stage1_col104[15] = fa_s0_c104_n766_s;
                stage1_col104[16] = fa_s0_c104_n767_s;
                stage1_col104[17] = fa_s0_c104_n768_s;
                stage1_col104[18] = fa_s0_c104_n769_s;
                stage1_col104[19] = fa_s0_c104_n770_s;
                stage1_col104[20] = fa_s0_c104_n771_s;
                stage1_col105[0] = fa_s0_c104_n761_c;
                stage1_col105[1] = fa_s0_c104_n762_c;
                stage1_col105[2] = fa_s0_c104_n763_c;
                stage1_col105[3] = fa_s0_c104_n764_c;
                stage1_col105[4] = fa_s0_c104_n765_c;
                stage1_col105[5] = fa_s0_c104_n766_c;
                stage1_col105[6] = fa_s0_c104_n767_c;
                stage1_col105[7] = fa_s0_c104_n768_c;
                stage1_col105[8] = fa_s0_c104_n769_c;
                stage1_col105[9] = fa_s0_c104_n770_c;
                stage1_col105[10] = fa_s0_c104_n771_c;
                stage1_col105[11] = fa_s0_c105_n772_s;
                stage1_col105[12] = fa_s0_c105_n773_s;
                stage1_col105[13] = fa_s0_c105_n774_s;
                stage1_col105[14] = fa_s0_c105_n775_s;
                stage1_col105[15] = fa_s0_c105_n776_s;
                stage1_col105[16] = fa_s0_c105_n777_s;
                stage1_col105[17] = fa_s0_c105_n778_s;
                stage1_col105[18] = fa_s0_c105_n779_s;
                stage1_col105[19] = fa_s0_c105_n780_s;
                stage1_col105[20] = fa_s0_c105_n781_s;
                stage1_col105[21] = stage0_col105[30];
                stage1_col105[22] = stage0_col105[31];
                stage1_col106[0] = fa_s0_c105_n772_c;
                stage1_col106[1] = fa_s0_c105_n773_c;
                stage1_col106[2] = fa_s0_c105_n774_c;
                stage1_col106[3] = fa_s0_c105_n775_c;
                stage1_col106[4] = fa_s0_c105_n776_c;
                stage1_col106[5] = fa_s0_c105_n777_c;
                stage1_col106[6] = fa_s0_c105_n778_c;
                stage1_col106[7] = fa_s0_c105_n779_c;
                stage1_col106[8] = fa_s0_c105_n780_c;
                stage1_col106[9] = fa_s0_c105_n781_c;
                stage1_col106[10] = fa_s0_c106_n782_s;
                stage1_col106[11] = fa_s0_c106_n783_s;
                stage1_col106[12] = fa_s0_c106_n784_s;
                stage1_col106[13] = fa_s0_c106_n785_s;
                stage1_col106[14] = fa_s0_c106_n786_s;
                stage1_col106[15] = fa_s0_c106_n787_s;
                stage1_col106[16] = fa_s0_c106_n788_s;
                stage1_col106[17] = fa_s0_c106_n789_s;
                stage1_col106[18] = fa_s0_c106_n790_s;
                stage1_col106[19] = fa_s0_c106_n791_s;
                stage1_col106[20] = fa_s0_c106_n792_s;
                stage1_col107[0] = fa_s0_c106_n782_c;
                stage1_col107[1] = fa_s0_c106_n783_c;
                stage1_col107[2] = fa_s0_c106_n784_c;
                stage1_col107[3] = fa_s0_c106_n785_c;
                stage1_col107[4] = fa_s0_c106_n786_c;
                stage1_col107[5] = fa_s0_c106_n787_c;
                stage1_col107[6] = fa_s0_c106_n788_c;
                stage1_col107[7] = fa_s0_c106_n789_c;
                stage1_col107[8] = fa_s0_c106_n790_c;
                stage1_col107[9] = fa_s0_c106_n791_c;
                stage1_col107[10] = fa_s0_c106_n792_c;
                stage1_col107[11] = fa_s0_c107_n793_s;
                stage1_col107[12] = fa_s0_c107_n794_s;
                stage1_col107[13] = fa_s0_c107_n795_s;
                stage1_col107[14] = fa_s0_c107_n796_s;
                stage1_col107[15] = fa_s0_c107_n797_s;
                stage1_col107[16] = fa_s0_c107_n798_s;
                stage1_col107[17] = fa_s0_c107_n799_s;
                stage1_col107[18] = fa_s0_c107_n800_s;
                stage1_col107[19] = fa_s0_c107_n801_s;
                stage1_col107[20] = fa_s0_c107_n802_s;
                stage1_col107[21] = stage0_col107[30];
                stage1_col107[22] = stage0_col107[31];
                stage1_col108[0] = fa_s0_c107_n793_c;
                stage1_col108[1] = fa_s0_c107_n794_c;
                stage1_col108[2] = fa_s0_c107_n795_c;
                stage1_col108[3] = fa_s0_c107_n796_c;
                stage1_col108[4] = fa_s0_c107_n797_c;
                stage1_col108[5] = fa_s0_c107_n798_c;
                stage1_col108[6] = fa_s0_c107_n799_c;
                stage1_col108[7] = fa_s0_c107_n800_c;
                stage1_col108[8] = fa_s0_c107_n801_c;
                stage1_col108[9] = fa_s0_c107_n802_c;
                stage1_col108[10] = fa_s0_c108_n803_s;
                stage1_col108[11] = fa_s0_c108_n804_s;
                stage1_col108[12] = fa_s0_c108_n805_s;
                stage1_col108[13] = fa_s0_c108_n806_s;
                stage1_col108[14] = fa_s0_c108_n807_s;
                stage1_col108[15] = fa_s0_c108_n808_s;
                stage1_col108[16] = fa_s0_c108_n809_s;
                stage1_col108[17] = fa_s0_c108_n810_s;
                stage1_col108[18] = fa_s0_c108_n811_s;
                stage1_col108[19] = fa_s0_c108_n812_s;
                stage1_col108[20] = fa_s0_c108_n813_s;
                stage1_col109[0] = fa_s0_c108_n803_c;
                stage1_col109[1] = fa_s0_c108_n804_c;
                stage1_col109[2] = fa_s0_c108_n805_c;
                stage1_col109[3] = fa_s0_c108_n806_c;
                stage1_col109[4] = fa_s0_c108_n807_c;
                stage1_col109[5] = fa_s0_c108_n808_c;
                stage1_col109[6] = fa_s0_c108_n809_c;
                stage1_col109[7] = fa_s0_c108_n810_c;
                stage1_col109[8] = fa_s0_c108_n811_c;
                stage1_col109[9] = fa_s0_c108_n812_c;
                stage1_col109[10] = fa_s0_c108_n813_c;
                stage1_col109[11] = fa_s0_c109_n814_s;
                stage1_col109[12] = fa_s0_c109_n815_s;
                stage1_col109[13] = fa_s0_c109_n816_s;
                stage1_col109[14] = fa_s0_c109_n817_s;
                stage1_col109[15] = fa_s0_c109_n818_s;
                stage1_col109[16] = fa_s0_c109_n819_s;
                stage1_col109[17] = fa_s0_c109_n820_s;
                stage1_col109[18] = fa_s0_c109_n821_s;
                stage1_col109[19] = fa_s0_c109_n822_s;
                stage1_col109[20] = fa_s0_c109_n823_s;
                stage1_col109[21] = stage0_col109[30];
                stage1_col109[22] = stage0_col109[31];
                stage1_col110[0] = fa_s0_c109_n814_c;
                stage1_col110[1] = fa_s0_c109_n815_c;
                stage1_col110[2] = fa_s0_c109_n816_c;
                stage1_col110[3] = fa_s0_c109_n817_c;
                stage1_col110[4] = fa_s0_c109_n818_c;
                stage1_col110[5] = fa_s0_c109_n819_c;
                stage1_col110[6] = fa_s0_c109_n820_c;
                stage1_col110[7] = fa_s0_c109_n821_c;
                stage1_col110[8] = fa_s0_c109_n822_c;
                stage1_col110[9] = fa_s0_c109_n823_c;
                stage1_col110[10] = fa_s0_c110_n824_s;
                stage1_col110[11] = fa_s0_c110_n825_s;
                stage1_col110[12] = fa_s0_c110_n826_s;
                stage1_col110[13] = fa_s0_c110_n827_s;
                stage1_col110[14] = fa_s0_c110_n828_s;
                stage1_col110[15] = fa_s0_c110_n829_s;
                stage1_col110[16] = fa_s0_c110_n830_s;
                stage1_col110[17] = fa_s0_c110_n831_s;
                stage1_col110[18] = fa_s0_c110_n832_s;
                stage1_col110[19] = fa_s0_c110_n833_s;
                stage1_col110[20] = fa_s0_c110_n834_s;
                stage1_col111[0] = fa_s0_c110_n824_c;
                stage1_col111[1] = fa_s0_c110_n825_c;
                stage1_col111[2] = fa_s0_c110_n826_c;
                stage1_col111[3] = fa_s0_c110_n827_c;
                stage1_col111[4] = fa_s0_c110_n828_c;
                stage1_col111[5] = fa_s0_c110_n829_c;
                stage1_col111[6] = fa_s0_c110_n830_c;
                stage1_col111[7] = fa_s0_c110_n831_c;
                stage1_col111[8] = fa_s0_c110_n832_c;
                stage1_col111[9] = fa_s0_c110_n833_c;
                stage1_col111[10] = fa_s0_c110_n834_c;
                stage1_col111[11] = fa_s0_c111_n835_s;
                stage1_col111[12] = fa_s0_c111_n836_s;
                stage1_col111[13] = fa_s0_c111_n837_s;
                stage1_col111[14] = fa_s0_c111_n838_s;
                stage1_col111[15] = fa_s0_c111_n839_s;
                stage1_col111[16] = fa_s0_c111_n840_s;
                stage1_col111[17] = fa_s0_c111_n841_s;
                stage1_col111[18] = fa_s0_c111_n842_s;
                stage1_col111[19] = fa_s0_c111_n843_s;
                stage1_col111[20] = fa_s0_c111_n844_s;
                stage1_col111[21] = stage0_col111[30];
                stage1_col111[22] = stage0_col111[31];
                stage1_col112[0] = fa_s0_c111_n835_c;
                stage1_col112[1] = fa_s0_c111_n836_c;
                stage1_col112[2] = fa_s0_c111_n837_c;
                stage1_col112[3] = fa_s0_c111_n838_c;
                stage1_col112[4] = fa_s0_c111_n839_c;
                stage1_col112[5] = fa_s0_c111_n840_c;
                stage1_col112[6] = fa_s0_c111_n841_c;
                stage1_col112[7] = fa_s0_c111_n842_c;
                stage1_col112[8] = fa_s0_c111_n843_c;
                stage1_col112[9] = fa_s0_c111_n844_c;
                stage1_col112[10] = fa_s0_c112_n845_s;
                stage1_col112[11] = fa_s0_c112_n846_s;
                stage1_col112[12] = fa_s0_c112_n847_s;
                stage1_col112[13] = fa_s0_c112_n848_s;
                stage1_col112[14] = fa_s0_c112_n849_s;
                stage1_col112[15] = fa_s0_c112_n850_s;
                stage1_col112[16] = fa_s0_c112_n851_s;
                stage1_col112[17] = fa_s0_c112_n852_s;
                stage1_col112[18] = fa_s0_c112_n853_s;
                stage1_col112[19] = fa_s0_c112_n854_s;
                stage1_col112[20] = fa_s0_c112_n855_s;
                stage1_col113[0] = fa_s0_c112_n845_c;
                stage1_col113[1] = fa_s0_c112_n846_c;
                stage1_col113[2] = fa_s0_c112_n847_c;
                stage1_col113[3] = fa_s0_c112_n848_c;
                stage1_col113[4] = fa_s0_c112_n849_c;
                stage1_col113[5] = fa_s0_c112_n850_c;
                stage1_col113[6] = fa_s0_c112_n851_c;
                stage1_col113[7] = fa_s0_c112_n852_c;
                stage1_col113[8] = fa_s0_c112_n853_c;
                stage1_col113[9] = fa_s0_c112_n854_c;
                stage1_col113[10] = fa_s0_c112_n855_c;
                stage1_col113[11] = fa_s0_c113_n856_s;
                stage1_col113[12] = fa_s0_c113_n857_s;
                stage1_col113[13] = fa_s0_c113_n858_s;
                stage1_col113[14] = fa_s0_c113_n859_s;
                stage1_col113[15] = fa_s0_c113_n860_s;
                stage1_col113[16] = fa_s0_c113_n861_s;
                stage1_col113[17] = fa_s0_c113_n862_s;
                stage1_col113[18] = fa_s0_c113_n863_s;
                stage1_col113[19] = fa_s0_c113_n864_s;
                stage1_col113[20] = fa_s0_c113_n865_s;
                stage1_col113[21] = stage0_col113[30];
                stage1_col113[22] = stage0_col113[31];
                stage1_col114[0] = fa_s0_c113_n856_c;
                stage1_col114[1] = fa_s0_c113_n857_c;
                stage1_col114[2] = fa_s0_c113_n858_c;
                stage1_col114[3] = fa_s0_c113_n859_c;
                stage1_col114[4] = fa_s0_c113_n860_c;
                stage1_col114[5] = fa_s0_c113_n861_c;
                stage1_col114[6] = fa_s0_c113_n862_c;
                stage1_col114[7] = fa_s0_c113_n863_c;
                stage1_col114[8] = fa_s0_c113_n864_c;
                stage1_col114[9] = fa_s0_c113_n865_c;
                stage1_col114[10] = fa_s0_c114_n866_s;
                stage1_col114[11] = fa_s0_c114_n867_s;
                stage1_col114[12] = fa_s0_c114_n868_s;
                stage1_col114[13] = fa_s0_c114_n869_s;
                stage1_col114[14] = fa_s0_c114_n870_s;
                stage1_col114[15] = fa_s0_c114_n871_s;
                stage1_col114[16] = fa_s0_c114_n872_s;
                stage1_col114[17] = fa_s0_c114_n873_s;
                stage1_col114[18] = fa_s0_c114_n874_s;
                stage1_col114[19] = fa_s0_c114_n875_s;
                stage1_col114[20] = fa_s0_c114_n876_s;
                stage1_col115[0] = fa_s0_c114_n866_c;
                stage1_col115[1] = fa_s0_c114_n867_c;
                stage1_col115[2] = fa_s0_c114_n868_c;
                stage1_col115[3] = fa_s0_c114_n869_c;
                stage1_col115[4] = fa_s0_c114_n870_c;
                stage1_col115[5] = fa_s0_c114_n871_c;
                stage1_col115[6] = fa_s0_c114_n872_c;
                stage1_col115[7] = fa_s0_c114_n873_c;
                stage1_col115[8] = fa_s0_c114_n874_c;
                stage1_col115[9] = fa_s0_c114_n875_c;
                stage1_col115[10] = fa_s0_c114_n876_c;
                stage1_col115[11] = fa_s0_c115_n877_s;
                stage1_col115[12] = fa_s0_c115_n878_s;
                stage1_col115[13] = fa_s0_c115_n879_s;
                stage1_col115[14] = fa_s0_c115_n880_s;
                stage1_col115[15] = fa_s0_c115_n881_s;
                stage1_col115[16] = fa_s0_c115_n882_s;
                stage1_col115[17] = fa_s0_c115_n883_s;
                stage1_col115[18] = fa_s0_c115_n884_s;
                stage1_col115[19] = fa_s0_c115_n885_s;
                stage1_col115[20] = fa_s0_c115_n886_s;
                stage1_col115[21] = stage0_col115[30];
                stage1_col115[22] = stage0_col115[31];
                stage1_col116[0] = fa_s0_c115_n877_c;
                stage1_col116[1] = fa_s0_c115_n878_c;
                stage1_col116[2] = fa_s0_c115_n879_c;
                stage1_col116[3] = fa_s0_c115_n880_c;
                stage1_col116[4] = fa_s0_c115_n881_c;
                stage1_col116[5] = fa_s0_c115_n882_c;
                stage1_col116[6] = fa_s0_c115_n883_c;
                stage1_col116[7] = fa_s0_c115_n884_c;
                stage1_col116[8] = fa_s0_c115_n885_c;
                stage1_col116[9] = fa_s0_c115_n886_c;
                stage1_col116[10] = fa_s0_c116_n887_s;
                stage1_col116[11] = fa_s0_c116_n888_s;
                stage1_col116[12] = fa_s0_c116_n889_s;
                stage1_col116[13] = fa_s0_c116_n890_s;
                stage1_col116[14] = fa_s0_c116_n891_s;
                stage1_col116[15] = fa_s0_c116_n892_s;
                stage1_col116[16] = fa_s0_c116_n893_s;
                stage1_col116[17] = fa_s0_c116_n894_s;
                stage1_col116[18] = fa_s0_c116_n895_s;
                stage1_col116[19] = fa_s0_c116_n896_s;
                stage1_col116[20] = fa_s0_c116_n897_s;
                stage1_col117[0] = fa_s0_c116_n887_c;
                stage1_col117[1] = fa_s0_c116_n888_c;
                stage1_col117[2] = fa_s0_c116_n889_c;
                stage1_col117[3] = fa_s0_c116_n890_c;
                stage1_col117[4] = fa_s0_c116_n891_c;
                stage1_col117[5] = fa_s0_c116_n892_c;
                stage1_col117[6] = fa_s0_c116_n893_c;
                stage1_col117[7] = fa_s0_c116_n894_c;
                stage1_col117[8] = fa_s0_c116_n895_c;
                stage1_col117[9] = fa_s0_c116_n896_c;
                stage1_col117[10] = fa_s0_c116_n897_c;
                stage1_col117[11] = fa_s0_c117_n898_s;
                stage1_col117[12] = fa_s0_c117_n899_s;
                stage1_col117[13] = fa_s0_c117_n900_s;
                stage1_col117[14] = fa_s0_c117_n901_s;
                stage1_col117[15] = fa_s0_c117_n902_s;
                stage1_col117[16] = fa_s0_c117_n903_s;
                stage1_col117[17] = fa_s0_c117_n904_s;
                stage1_col117[18] = fa_s0_c117_n905_s;
                stage1_col117[19] = fa_s0_c117_n906_s;
                stage1_col117[20] = fa_s0_c117_n907_s;
                stage1_col117[21] = stage0_col117[30];
                stage1_col117[22] = stage0_col117[31];
                stage1_col118[0] = fa_s0_c117_n898_c;
                stage1_col118[1] = fa_s0_c117_n899_c;
                stage1_col118[2] = fa_s0_c117_n900_c;
                stage1_col118[3] = fa_s0_c117_n901_c;
                stage1_col118[4] = fa_s0_c117_n902_c;
                stage1_col118[5] = fa_s0_c117_n903_c;
                stage1_col118[6] = fa_s0_c117_n904_c;
                stage1_col118[7] = fa_s0_c117_n905_c;
                stage1_col118[8] = fa_s0_c117_n906_c;
                stage1_col118[9] = fa_s0_c117_n907_c;
                stage1_col118[10] = fa_s0_c118_n908_s;
                stage1_col118[11] = fa_s0_c118_n909_s;
                stage1_col118[12] = fa_s0_c118_n910_s;
                stage1_col118[13] = fa_s0_c118_n911_s;
                stage1_col118[14] = fa_s0_c118_n912_s;
                stage1_col118[15] = fa_s0_c118_n913_s;
                stage1_col118[16] = fa_s0_c118_n914_s;
                stage1_col118[17] = fa_s0_c118_n915_s;
                stage1_col118[18] = fa_s0_c118_n916_s;
                stage1_col118[19] = fa_s0_c118_n917_s;
                stage1_col118[20] = fa_s0_c118_n918_s;
                stage1_col119[0] = fa_s0_c118_n908_c;
                stage1_col119[1] = fa_s0_c118_n909_c;
                stage1_col119[2] = fa_s0_c118_n910_c;
                stage1_col119[3] = fa_s0_c118_n911_c;
                stage1_col119[4] = fa_s0_c118_n912_c;
                stage1_col119[5] = fa_s0_c118_n913_c;
                stage1_col119[6] = fa_s0_c118_n914_c;
                stage1_col119[7] = fa_s0_c118_n915_c;
                stage1_col119[8] = fa_s0_c118_n916_c;
                stage1_col119[9] = fa_s0_c118_n917_c;
                stage1_col119[10] = fa_s0_c118_n918_c;
                stage1_col119[11] = fa_s0_c119_n919_s;
                stage1_col119[12] = fa_s0_c119_n920_s;
                stage1_col119[13] = fa_s0_c119_n921_s;
                stage1_col119[14] = fa_s0_c119_n922_s;
                stage1_col119[15] = fa_s0_c119_n923_s;
                stage1_col119[16] = fa_s0_c119_n924_s;
                stage1_col119[17] = fa_s0_c119_n925_s;
                stage1_col119[18] = fa_s0_c119_n926_s;
                stage1_col119[19] = fa_s0_c119_n927_s;
                stage1_col119[20] = fa_s0_c119_n928_s;
                stage1_col119[21] = stage0_col119[30];
                stage1_col119[22] = stage0_col119[31];
                stage1_col120[0] = fa_s0_c119_n919_c;
                stage1_col120[1] = fa_s0_c119_n920_c;
                stage1_col120[2] = fa_s0_c119_n921_c;
                stage1_col120[3] = fa_s0_c119_n922_c;
                stage1_col120[4] = fa_s0_c119_n923_c;
                stage1_col120[5] = fa_s0_c119_n924_c;
                stage1_col120[6] = fa_s0_c119_n925_c;
                stage1_col120[7] = fa_s0_c119_n926_c;
                stage1_col120[8] = fa_s0_c119_n927_c;
                stage1_col120[9] = fa_s0_c119_n928_c;
                stage1_col120[10] = fa_s0_c120_n929_s;
                stage1_col120[11] = fa_s0_c120_n930_s;
                stage1_col120[12] = fa_s0_c120_n931_s;
                stage1_col120[13] = fa_s0_c120_n932_s;
                stage1_col120[14] = fa_s0_c120_n933_s;
                stage1_col120[15] = fa_s0_c120_n934_s;
                stage1_col120[16] = fa_s0_c120_n935_s;
                stage1_col120[17] = fa_s0_c120_n936_s;
                stage1_col120[18] = fa_s0_c120_n937_s;
                stage1_col120[19] = fa_s0_c120_n938_s;
                stage1_col120[20] = fa_s0_c120_n939_s;
                stage1_col121[0] = fa_s0_c120_n929_c;
                stage1_col121[1] = fa_s0_c120_n930_c;
                stage1_col121[2] = fa_s0_c120_n931_c;
                stage1_col121[3] = fa_s0_c120_n932_c;
                stage1_col121[4] = fa_s0_c120_n933_c;
                stage1_col121[5] = fa_s0_c120_n934_c;
                stage1_col121[6] = fa_s0_c120_n935_c;
                stage1_col121[7] = fa_s0_c120_n936_c;
                stage1_col121[8] = fa_s0_c120_n937_c;
                stage1_col121[9] = fa_s0_c120_n938_c;
                stage1_col121[10] = fa_s0_c120_n939_c;
                stage1_col121[11] = fa_s0_c121_n940_s;
                stage1_col121[12] = fa_s0_c121_n941_s;
                stage1_col121[13] = fa_s0_c121_n942_s;
                stage1_col121[14] = fa_s0_c121_n943_s;
                stage1_col121[15] = fa_s0_c121_n944_s;
                stage1_col121[16] = fa_s0_c121_n945_s;
                stage1_col121[17] = fa_s0_c121_n946_s;
                stage1_col121[18] = fa_s0_c121_n947_s;
                stage1_col121[19] = fa_s0_c121_n948_s;
                stage1_col121[20] = fa_s0_c121_n949_s;
                stage1_col121[21] = stage0_col121[30];
                stage1_col121[22] = stage0_col121[31];
                stage1_col122[0] = fa_s0_c121_n940_c;
                stage1_col122[1] = fa_s0_c121_n941_c;
                stage1_col122[2] = fa_s0_c121_n942_c;
                stage1_col122[3] = fa_s0_c121_n943_c;
                stage1_col122[4] = fa_s0_c121_n944_c;
                stage1_col122[5] = fa_s0_c121_n945_c;
                stage1_col122[6] = fa_s0_c121_n946_c;
                stage1_col122[7] = fa_s0_c121_n947_c;
                stage1_col122[8] = fa_s0_c121_n948_c;
                stage1_col122[9] = fa_s0_c121_n949_c;
                stage1_col122[10] = fa_s0_c122_n950_s;
                stage1_col122[11] = fa_s0_c122_n951_s;
                stage1_col122[12] = fa_s0_c122_n952_s;
                stage1_col122[13] = fa_s0_c122_n953_s;
                stage1_col122[14] = fa_s0_c122_n954_s;
                stage1_col122[15] = fa_s0_c122_n955_s;
                stage1_col122[16] = fa_s0_c122_n956_s;
                stage1_col122[17] = fa_s0_c122_n957_s;
                stage1_col122[18] = fa_s0_c122_n958_s;
                stage1_col122[19] = fa_s0_c122_n959_s;
                stage1_col122[20] = fa_s0_c122_n960_s;
                stage1_col123[0] = fa_s0_c122_n950_c;
                stage1_col123[1] = fa_s0_c122_n951_c;
                stage1_col123[2] = fa_s0_c122_n952_c;
                stage1_col123[3] = fa_s0_c122_n953_c;
                stage1_col123[4] = fa_s0_c122_n954_c;
                stage1_col123[5] = fa_s0_c122_n955_c;
                stage1_col123[6] = fa_s0_c122_n956_c;
                stage1_col123[7] = fa_s0_c122_n957_c;
                stage1_col123[8] = fa_s0_c122_n958_c;
                stage1_col123[9] = fa_s0_c122_n959_c;
                stage1_col123[10] = fa_s0_c122_n960_c;
                stage1_col123[11] = fa_s0_c123_n961_s;
                stage1_col123[12] = fa_s0_c123_n962_s;
                stage1_col123[13] = fa_s0_c123_n963_s;
                stage1_col123[14] = fa_s0_c123_n964_s;
                stage1_col123[15] = fa_s0_c123_n965_s;
                stage1_col123[16] = fa_s0_c123_n966_s;
                stage1_col123[17] = fa_s0_c123_n967_s;
                stage1_col123[18] = fa_s0_c123_n968_s;
                stage1_col123[19] = fa_s0_c123_n969_s;
                stage1_col123[20] = fa_s0_c123_n970_s;
                stage1_col123[21] = stage0_col123[30];
                stage1_col123[22] = stage0_col123[31];
                stage1_col124[0] = fa_s0_c123_n961_c;
                stage1_col124[1] = fa_s0_c123_n962_c;
                stage1_col124[2] = fa_s0_c123_n963_c;
                stage1_col124[3] = fa_s0_c123_n964_c;
                stage1_col124[4] = fa_s0_c123_n965_c;
                stage1_col124[5] = fa_s0_c123_n966_c;
                stage1_col124[6] = fa_s0_c123_n967_c;
                stage1_col124[7] = fa_s0_c123_n968_c;
                stage1_col124[8] = fa_s0_c123_n969_c;
                stage1_col124[9] = fa_s0_c123_n970_c;
                stage1_col124[10] = fa_s0_c124_n971_s;
                stage1_col124[11] = fa_s0_c124_n972_s;
                stage1_col124[12] = fa_s0_c124_n973_s;
                stage1_col124[13] = fa_s0_c124_n974_s;
                stage1_col124[14] = fa_s0_c124_n975_s;
                stage1_col124[15] = fa_s0_c124_n976_s;
                stage1_col124[16] = fa_s0_c124_n977_s;
                stage1_col124[17] = fa_s0_c124_n978_s;
                stage1_col124[18] = fa_s0_c124_n979_s;
                stage1_col124[19] = fa_s0_c124_n980_s;
                stage1_col124[20] = fa_s0_c124_n981_s;
                stage1_col125[0] = fa_s0_c124_n971_c;
                stage1_col125[1] = fa_s0_c124_n972_c;
                stage1_col125[2] = fa_s0_c124_n973_c;
                stage1_col125[3] = fa_s0_c124_n974_c;
                stage1_col125[4] = fa_s0_c124_n975_c;
                stage1_col125[5] = fa_s0_c124_n976_c;
                stage1_col125[6] = fa_s0_c124_n977_c;
                stage1_col125[7] = fa_s0_c124_n978_c;
                stage1_col125[8] = fa_s0_c124_n979_c;
                stage1_col125[9] = fa_s0_c124_n980_c;
                stage1_col125[10] = fa_s0_c124_n981_c;
                stage1_col125[11] = fa_s0_c125_n982_s;
                stage1_col125[12] = fa_s0_c125_n983_s;
                stage1_col125[13] = fa_s0_c125_n984_s;
                stage1_col125[14] = fa_s0_c125_n985_s;
                stage1_col125[15] = fa_s0_c125_n986_s;
                stage1_col125[16] = fa_s0_c125_n987_s;
                stage1_col125[17] = fa_s0_c125_n988_s;
                stage1_col125[18] = fa_s0_c125_n989_s;
                stage1_col125[19] = fa_s0_c125_n990_s;
                stage1_col125[20] = fa_s0_c125_n991_s;
                stage1_col125[21] = stage0_col125[0];
                stage1_col125[22] = stage0_col125[31];
                stage1_col126[0] = fa_s0_c125_n982_c;
                stage1_col126[1] = fa_s0_c125_n983_c;
                stage1_col126[2] = fa_s0_c125_n984_c;
                stage1_col126[3] = fa_s0_c125_n985_c;
                stage1_col126[4] = fa_s0_c125_n986_c;
                stage1_col126[5] = fa_s0_c125_n987_c;
                stage1_col126[6] = fa_s0_c125_n988_c;
                stage1_col126[7] = fa_s0_c125_n989_c;
                stage1_col126[8] = fa_s0_c125_n990_c;
                stage1_col126[9] = fa_s0_c125_n991_c;
                stage1_col126[10] = fa_s0_c126_n992_s;
                stage1_col126[11] = fa_s0_c126_n993_s;
                stage1_col126[12] = fa_s0_c126_n994_s;
                stage1_col126[13] = fa_s0_c126_n995_s;
                stage1_col126[14] = fa_s0_c126_n996_s;
                stage1_col126[15] = fa_s0_c126_n997_s;
                stage1_col126[16] = fa_s0_c126_n998_s;
                stage1_col126[17] = fa_s0_c126_n999_s;
                stage1_col126[18] = fa_s0_c126_n1000_s;
                stage1_col126[19] = fa_s0_c126_n1001_s;
                stage1_col126[20] = fa_s0_c126_n1002_s;
                stage1_col127[0] = fa_s0_c126_n992_c;
                stage1_col127[1] = fa_s0_c126_n993_c;
                stage1_col127[2] = fa_s0_c126_n994_c;
                stage1_col127[3] = fa_s0_c126_n995_c;
                stage1_col127[4] = fa_s0_c126_n996_c;
                stage1_col127[5] = fa_s0_c126_n997_c;
                stage1_col127[6] = fa_s0_c126_n998_c;
                stage1_col127[7] = fa_s0_c126_n999_c;
                stage1_col127[8] = fa_s0_c126_n1000_c;
                stage1_col127[9] = fa_s0_c126_n1001_c;
                stage1_col127[10] = fa_s0_c126_n1002_c;
                stage1_col127[11] = stage0_col127[0];
                stage1_col127[12] = stage0_col127[0];
                stage1_col127[13] = stage0_col127[0];
                stage1_col127[14] = stage0_col127[0];
                stage1_col127[15] = stage0_col127[0];
                stage1_col127[16] = stage0_col127[0];
                stage1_col127[17] = stage0_col127[0];
                stage1_col127[18] = stage0_col127[0];
                stage1_col127[19] = stage0_col127[0];
                stage1_col127[20] = stage0_col127[0];
                stage1_col127[21] = stage0_col127[0];
                stage1_col127[22] = stage0_col127[0];
                stage1_col127[23] = stage0_col127[0];
                stage1_col127[24] = stage0_col127[0];
                stage1_col127[25] = stage0_col127[0];
                stage1_col127[26] = stage0_col127[0];
                stage1_col127[27] = stage0_col127[0];
                stage1_col127[28] = stage0_col127[0];
                stage1_col127[29] = stage0_col127[0];
                stage1_col127[30] = stage0_col127[0];
                stage1_col127[31] = stage0_col127[0];
                stage1_col127[32] = stage0_col127[0];
                stage1_col127[33] = stage0_col127[0];
                stage1_col127[34] = stage0_col127[0];
                stage1_col127[35] = stage0_col127[0];
                stage1_col127[36] = stage0_col127[0];
                stage1_col127[37] = stage0_col127[0];
                stage1_col127[38] = stage0_col127[0];
                stage1_col127[39] = stage0_col127[0];
                stage1_col127[40] = stage0_col127[0];
                stage1_col127[41] = stage0_col127[0];
                stage1_col127[42] = stage0_col127[0];
            end
        end
    endgenerate

    // Stage 2: Reduction
    fa fa_s1_c3_n0 (
        .a(stage1_col3[0]),
        .b(stage1_col3[1]),
        .c_in(stage1_col3[2]),
        .s(fa_s1_c3_n0_s),
        .c_out(fa_s1_c3_n0_c)
    );

    fa fa_s1_c6_n1 (
        .a(stage1_col6[0]),
        .b(stage1_col6[1]),
        .c_in(stage1_col6[2]),
        .s(fa_s1_c6_n1_s),
        .c_out(fa_s1_c6_n1_c)
    );

    fa fa_s1_c7_n2 (
        .a(stage1_col7[0]),
        .b(stage1_col7[1]),
        .c_in(stage1_col7[2]),
        .s(fa_s1_c7_n2_s),
        .c_out(fa_s1_c7_n2_c)
    );

    fa fa_s1_c8_n3 (
        .a(stage1_col8[0]),
        .b(stage1_col8[1]),
        .c_in(stage1_col8[2]),
        .s(fa_s1_c8_n3_s),
        .c_out(fa_s1_c8_n3_c)
    );

    fa fa_s1_c9_n4 (
        .a(stage1_col9[0]),
        .b(stage1_col9[1]),
        .c_in(stage1_col9[2]),
        .s(fa_s1_c9_n4_s),
        .c_out(fa_s1_c9_n4_c)
    );

    fa fa_s1_c10_n5 (
        .a(stage1_col10[0]),
        .b(stage1_col10[1]),
        .c_in(stage1_col10[2]),
        .s(fa_s1_c10_n5_s),
        .c_out(fa_s1_c10_n5_c)
    );

    fa fa_s1_c11_n6 (
        .a(stage1_col11[0]),
        .b(stage1_col11[1]),
        .c_in(stage1_col11[2]),
        .s(fa_s1_c11_n6_s),
        .c_out(fa_s1_c11_n6_c)
    );

    fa fa_s1_c12_n7 (
        .a(stage1_col12[0]),
        .b(stage1_col12[1]),
        .c_in(stage1_col12[2]),
        .s(fa_s1_c12_n7_s),
        .c_out(fa_s1_c12_n7_c)
    );

    fa fa_s1_c12_n8 (
        .a(stage1_col12[3]),
        .b(stage1_col12[4]),
        .c_in(stage1_col12[5]),
        .s(fa_s1_c12_n8_s),
        .c_out(fa_s1_c12_n8_c)
    );

    fa fa_s1_c13_n9 (
        .a(stage1_col13[0]),
        .b(stage1_col13[1]),
        .c_in(stage1_col13[2]),
        .s(fa_s1_c13_n9_s),
        .c_out(fa_s1_c13_n9_c)
    );

    fa fa_s1_c14_n10 (
        .a(stage1_col14[0]),
        .b(stage1_col14[1]),
        .c_in(stage1_col14[2]),
        .s(fa_s1_c14_n10_s),
        .c_out(fa_s1_c14_n10_c)
    );

    fa fa_s1_c15_n11 (
        .a(stage1_col15[0]),
        .b(stage1_col15[1]),
        .c_in(stage1_col15[2]),
        .s(fa_s1_c15_n11_s),
        .c_out(fa_s1_c15_n11_c)
    );

    fa fa_s1_c15_n12 (
        .a(stage1_col15[3]),
        .b(stage1_col15[4]),
        .c_in(stage1_col15[5]),
        .s(fa_s1_c15_n12_s),
        .c_out(fa_s1_c15_n12_c)
    );

    fa fa_s1_c16_n13 (
        .a(stage1_col16[0]),
        .b(stage1_col16[1]),
        .c_in(stage1_col16[2]),
        .s(fa_s1_c16_n13_s),
        .c_out(fa_s1_c16_n13_c)
    );

    fa fa_s1_c16_n14 (
        .a(stage1_col16[3]),
        .b(stage1_col16[4]),
        .c_in(stage1_col16[5]),
        .s(fa_s1_c16_n14_s),
        .c_out(fa_s1_c16_n14_c)
    );

    fa fa_s1_c17_n15 (
        .a(stage1_col17[0]),
        .b(stage1_col17[1]),
        .c_in(stage1_col17[2]),
        .s(fa_s1_c17_n15_s),
        .c_out(fa_s1_c17_n15_c)
    );

    fa fa_s1_c17_n16 (
        .a(stage1_col17[3]),
        .b(stage1_col17[4]),
        .c_in(stage1_col17[5]),
        .s(fa_s1_c17_n16_s),
        .c_out(fa_s1_c17_n16_c)
    );

    fa fa_s1_c18_n17 (
        .a(stage1_col18[0]),
        .b(stage1_col18[1]),
        .c_in(stage1_col18[2]),
        .s(fa_s1_c18_n17_s),
        .c_out(fa_s1_c18_n17_c)
    );

    fa fa_s1_c18_n18 (
        .a(stage1_col18[3]),
        .b(stage1_col18[4]),
        .c_in(stage1_col18[5]),
        .s(fa_s1_c18_n18_s),
        .c_out(fa_s1_c18_n18_c)
    );

    fa fa_s1_c19_n19 (
        .a(stage1_col19[0]),
        .b(stage1_col19[1]),
        .c_in(stage1_col19[2]),
        .s(fa_s1_c19_n19_s),
        .c_out(fa_s1_c19_n19_c)
    );

    fa fa_s1_c19_n20 (
        .a(stage1_col19[3]),
        .b(stage1_col19[4]),
        .c_in(stage1_col19[5]),
        .s(fa_s1_c19_n20_s),
        .c_out(fa_s1_c19_n20_c)
    );

    fa fa_s1_c20_n21 (
        .a(stage1_col20[0]),
        .b(stage1_col20[1]),
        .c_in(stage1_col20[2]),
        .s(fa_s1_c20_n21_s),
        .c_out(fa_s1_c20_n21_c)
    );

    fa fa_s1_c20_n22 (
        .a(stage1_col20[3]),
        .b(stage1_col20[4]),
        .c_in(stage1_col20[5]),
        .s(fa_s1_c20_n22_s),
        .c_out(fa_s1_c20_n22_c)
    );

    fa fa_s1_c21_n23 (
        .a(stage1_col21[0]),
        .b(stage1_col21[1]),
        .c_in(stage1_col21[2]),
        .s(fa_s1_c21_n23_s),
        .c_out(fa_s1_c21_n23_c)
    );

    fa fa_s1_c21_n24 (
        .a(stage1_col21[3]),
        .b(stage1_col21[4]),
        .c_in(stage1_col21[5]),
        .s(fa_s1_c21_n24_s),
        .c_out(fa_s1_c21_n24_c)
    );

    fa fa_s1_c21_n25 (
        .a(stage1_col21[6]),
        .b(stage1_col21[7]),
        .c_in(stage1_col21[8]),
        .s(fa_s1_c21_n25_s),
        .c_out(fa_s1_c21_n25_c)
    );

    fa fa_s1_c22_n26 (
        .a(stage1_col22[0]),
        .b(stage1_col22[1]),
        .c_in(stage1_col22[2]),
        .s(fa_s1_c22_n26_s),
        .c_out(fa_s1_c22_n26_c)
    );

    fa fa_s1_c22_n27 (
        .a(stage1_col22[3]),
        .b(stage1_col22[4]),
        .c_in(stage1_col22[5]),
        .s(fa_s1_c22_n27_s),
        .c_out(fa_s1_c22_n27_c)
    );

    fa fa_s1_c23_n28 (
        .a(stage1_col23[0]),
        .b(stage1_col23[1]),
        .c_in(stage1_col23[2]),
        .s(fa_s1_c23_n28_s),
        .c_out(fa_s1_c23_n28_c)
    );

    fa fa_s1_c23_n29 (
        .a(stage1_col23[3]),
        .b(stage1_col23[4]),
        .c_in(stage1_col23[5]),
        .s(fa_s1_c23_n29_s),
        .c_out(fa_s1_c23_n29_c)
    );

    fa fa_s1_c24_n30 (
        .a(stage1_col24[0]),
        .b(stage1_col24[1]),
        .c_in(stage1_col24[2]),
        .s(fa_s1_c24_n30_s),
        .c_out(fa_s1_c24_n30_c)
    );

    fa fa_s1_c24_n31 (
        .a(stage1_col24[3]),
        .b(stage1_col24[4]),
        .c_in(stage1_col24[5]),
        .s(fa_s1_c24_n31_s),
        .c_out(fa_s1_c24_n31_c)
    );

    fa fa_s1_c24_n32 (
        .a(stage1_col24[6]),
        .b(stage1_col24[7]),
        .c_in(stage1_col24[8]),
        .s(fa_s1_c24_n32_s),
        .c_out(fa_s1_c24_n32_c)
    );

    fa fa_s1_c25_n33 (
        .a(stage1_col25[0]),
        .b(stage1_col25[1]),
        .c_in(stage1_col25[2]),
        .s(fa_s1_c25_n33_s),
        .c_out(fa_s1_c25_n33_c)
    );

    fa fa_s1_c25_n34 (
        .a(stage1_col25[3]),
        .b(stage1_col25[4]),
        .c_in(stage1_col25[5]),
        .s(fa_s1_c25_n34_s),
        .c_out(fa_s1_c25_n34_c)
    );

    fa fa_s1_c25_n35 (
        .a(stage1_col25[6]),
        .b(stage1_col25[7]),
        .c_in(stage1_col25[8]),
        .s(fa_s1_c25_n35_s),
        .c_out(fa_s1_c25_n35_c)
    );

    fa fa_s1_c26_n36 (
        .a(stage1_col26[0]),
        .b(stage1_col26[1]),
        .c_in(stage1_col26[2]),
        .s(fa_s1_c26_n36_s),
        .c_out(fa_s1_c26_n36_c)
    );

    fa fa_s1_c26_n37 (
        .a(stage1_col26[3]),
        .b(stage1_col26[4]),
        .c_in(stage1_col26[5]),
        .s(fa_s1_c26_n37_s),
        .c_out(fa_s1_c26_n37_c)
    );

    fa fa_s1_c26_n38 (
        .a(stage1_col26[6]),
        .b(stage1_col26[7]),
        .c_in(stage1_col26[8]),
        .s(fa_s1_c26_n38_s),
        .c_out(fa_s1_c26_n38_c)
    );

    fa fa_s1_c27_n39 (
        .a(stage1_col27[0]),
        .b(stage1_col27[1]),
        .c_in(stage1_col27[2]),
        .s(fa_s1_c27_n39_s),
        .c_out(fa_s1_c27_n39_c)
    );

    fa fa_s1_c27_n40 (
        .a(stage1_col27[3]),
        .b(stage1_col27[4]),
        .c_in(stage1_col27[5]),
        .s(fa_s1_c27_n40_s),
        .c_out(fa_s1_c27_n40_c)
    );

    fa fa_s1_c27_n41 (
        .a(stage1_col27[6]),
        .b(stage1_col27[7]),
        .c_in(stage1_col27[8]),
        .s(fa_s1_c27_n41_s),
        .c_out(fa_s1_c27_n41_c)
    );

    fa fa_s1_c28_n42 (
        .a(stage1_col28[0]),
        .b(stage1_col28[1]),
        .c_in(stage1_col28[2]),
        .s(fa_s1_c28_n42_s),
        .c_out(fa_s1_c28_n42_c)
    );

    fa fa_s1_c28_n43 (
        .a(stage1_col28[3]),
        .b(stage1_col28[4]),
        .c_in(stage1_col28[5]),
        .s(fa_s1_c28_n43_s),
        .c_out(fa_s1_c28_n43_c)
    );

    fa fa_s1_c28_n44 (
        .a(stage1_col28[6]),
        .b(stage1_col28[7]),
        .c_in(stage1_col28[8]),
        .s(fa_s1_c28_n44_s),
        .c_out(fa_s1_c28_n44_c)
    );

    fa fa_s1_c29_n45 (
        .a(stage1_col29[0]),
        .b(stage1_col29[1]),
        .c_in(stage1_col29[2]),
        .s(fa_s1_c29_n45_s),
        .c_out(fa_s1_c29_n45_c)
    );

    fa fa_s1_c29_n46 (
        .a(stage1_col29[3]),
        .b(stage1_col29[4]),
        .c_in(stage1_col29[5]),
        .s(fa_s1_c29_n46_s),
        .c_out(fa_s1_c29_n46_c)
    );

    fa fa_s1_c29_n47 (
        .a(stage1_col29[6]),
        .b(stage1_col29[7]),
        .c_in(stage1_col29[8]),
        .s(fa_s1_c29_n47_s),
        .c_out(fa_s1_c29_n47_c)
    );

    fa fa_s1_c30_n48 (
        .a(stage1_col30[0]),
        .b(stage1_col30[1]),
        .c_in(stage1_col30[2]),
        .s(fa_s1_c30_n48_s),
        .c_out(fa_s1_c30_n48_c)
    );

    fa fa_s1_c30_n49 (
        .a(stage1_col30[3]),
        .b(stage1_col30[4]),
        .c_in(stage1_col30[5]),
        .s(fa_s1_c30_n49_s),
        .c_out(fa_s1_c30_n49_c)
    );

    fa fa_s1_c30_n50 (
        .a(stage1_col30[6]),
        .b(stage1_col30[7]),
        .c_in(stage1_col30[8]),
        .s(fa_s1_c30_n50_s),
        .c_out(fa_s1_c30_n50_c)
    );

    fa fa_s1_c30_n51 (
        .a(stage1_col30[9]),
        .b(stage1_col30[10]),
        .c_in(stage1_col30[11]),
        .s(fa_s1_c30_n51_s),
        .c_out(fa_s1_c30_n51_c)
    );

    fa fa_s1_c31_n52 (
        .a(stage1_col31[0]),
        .b(stage1_col31[1]),
        .c_in(stage1_col31[2]),
        .s(fa_s1_c31_n52_s),
        .c_out(fa_s1_c31_n52_c)
    );

    fa fa_s1_c31_n53 (
        .a(stage1_col31[3]),
        .b(stage1_col31[4]),
        .c_in(stage1_col31[5]),
        .s(fa_s1_c31_n53_s),
        .c_out(fa_s1_c31_n53_c)
    );

    fa fa_s1_c31_n54 (
        .a(stage1_col31[6]),
        .b(stage1_col31[7]),
        .c_in(stage1_col31[8]),
        .s(fa_s1_c31_n54_s),
        .c_out(fa_s1_c31_n54_c)
    );

    fa fa_s1_c32_n55 (
        .a(stage1_col32[0]),
        .b(stage1_col32[1]),
        .c_in(stage1_col32[2]),
        .s(fa_s1_c32_n55_s),
        .c_out(fa_s1_c32_n55_c)
    );

    fa fa_s1_c32_n56 (
        .a(stage1_col32[3]),
        .b(stage1_col32[4]),
        .c_in(stage1_col32[5]),
        .s(fa_s1_c32_n56_s),
        .c_out(fa_s1_c32_n56_c)
    );

    fa fa_s1_c32_n57 (
        .a(stage1_col32[6]),
        .b(stage1_col32[7]),
        .c_in(stage1_col32[8]),
        .s(fa_s1_c32_n57_s),
        .c_out(fa_s1_c32_n57_c)
    );

    fa fa_s1_c33_n58 (
        .a(stage1_col33[0]),
        .b(stage1_col33[1]),
        .c_in(stage1_col33[2]),
        .s(fa_s1_c33_n58_s),
        .c_out(fa_s1_c33_n58_c)
    );

    fa fa_s1_c33_n59 (
        .a(stage1_col33[3]),
        .b(stage1_col33[4]),
        .c_in(stage1_col33[5]),
        .s(fa_s1_c33_n59_s),
        .c_out(fa_s1_c33_n59_c)
    );

    fa fa_s1_c33_n60 (
        .a(stage1_col33[6]),
        .b(stage1_col33[7]),
        .c_in(stage1_col33[8]),
        .s(fa_s1_c33_n60_s),
        .c_out(fa_s1_c33_n60_c)
    );

    fa fa_s1_c33_n61 (
        .a(stage1_col33[9]),
        .b(stage1_col33[10]),
        .c_in(stage1_col33[11]),
        .s(fa_s1_c33_n61_s),
        .c_out(fa_s1_c33_n61_c)
    );

    fa fa_s1_c34_n62 (
        .a(stage1_col34[0]),
        .b(stage1_col34[1]),
        .c_in(stage1_col34[2]),
        .s(fa_s1_c34_n62_s),
        .c_out(fa_s1_c34_n62_c)
    );

    fa fa_s1_c34_n63 (
        .a(stage1_col34[3]),
        .b(stage1_col34[4]),
        .c_in(stage1_col34[5]),
        .s(fa_s1_c34_n63_s),
        .c_out(fa_s1_c34_n63_c)
    );

    fa fa_s1_c34_n64 (
        .a(stage1_col34[6]),
        .b(stage1_col34[7]),
        .c_in(stage1_col34[8]),
        .s(fa_s1_c34_n64_s),
        .c_out(fa_s1_c34_n64_c)
    );

    fa fa_s1_c34_n65 (
        .a(stage1_col34[9]),
        .b(stage1_col34[10]),
        .c_in(stage1_col34[11]),
        .s(fa_s1_c34_n65_s),
        .c_out(fa_s1_c34_n65_c)
    );

    fa fa_s1_c35_n66 (
        .a(stage1_col35[0]),
        .b(stage1_col35[1]),
        .c_in(stage1_col35[2]),
        .s(fa_s1_c35_n66_s),
        .c_out(fa_s1_c35_n66_c)
    );

    fa fa_s1_c35_n67 (
        .a(stage1_col35[3]),
        .b(stage1_col35[4]),
        .c_in(stage1_col35[5]),
        .s(fa_s1_c35_n67_s),
        .c_out(fa_s1_c35_n67_c)
    );

    fa fa_s1_c35_n68 (
        .a(stage1_col35[6]),
        .b(stage1_col35[7]),
        .c_in(stage1_col35[8]),
        .s(fa_s1_c35_n68_s),
        .c_out(fa_s1_c35_n68_c)
    );

    fa fa_s1_c35_n69 (
        .a(stage1_col35[9]),
        .b(stage1_col35[10]),
        .c_in(stage1_col35[11]),
        .s(fa_s1_c35_n69_s),
        .c_out(fa_s1_c35_n69_c)
    );

    fa fa_s1_c36_n70 (
        .a(stage1_col36[0]),
        .b(stage1_col36[1]),
        .c_in(stage1_col36[2]),
        .s(fa_s1_c36_n70_s),
        .c_out(fa_s1_c36_n70_c)
    );

    fa fa_s1_c36_n71 (
        .a(stage1_col36[3]),
        .b(stage1_col36[4]),
        .c_in(stage1_col36[5]),
        .s(fa_s1_c36_n71_s),
        .c_out(fa_s1_c36_n71_c)
    );

    fa fa_s1_c36_n72 (
        .a(stage1_col36[6]),
        .b(stage1_col36[7]),
        .c_in(stage1_col36[8]),
        .s(fa_s1_c36_n72_s),
        .c_out(fa_s1_c36_n72_c)
    );

    fa fa_s1_c36_n73 (
        .a(stage1_col36[9]),
        .b(stage1_col36[10]),
        .c_in(stage1_col36[11]),
        .s(fa_s1_c36_n73_s),
        .c_out(fa_s1_c36_n73_c)
    );

    fa fa_s1_c37_n74 (
        .a(stage1_col37[0]),
        .b(stage1_col37[1]),
        .c_in(stage1_col37[2]),
        .s(fa_s1_c37_n74_s),
        .c_out(fa_s1_c37_n74_c)
    );

    fa fa_s1_c37_n75 (
        .a(stage1_col37[3]),
        .b(stage1_col37[4]),
        .c_in(stage1_col37[5]),
        .s(fa_s1_c37_n75_s),
        .c_out(fa_s1_c37_n75_c)
    );

    fa fa_s1_c37_n76 (
        .a(stage1_col37[6]),
        .b(stage1_col37[7]),
        .c_in(stage1_col37[8]),
        .s(fa_s1_c37_n76_s),
        .c_out(fa_s1_c37_n76_c)
    );

    fa fa_s1_c37_n77 (
        .a(stage1_col37[9]),
        .b(stage1_col37[10]),
        .c_in(stage1_col37[11]),
        .s(fa_s1_c37_n77_s),
        .c_out(fa_s1_c37_n77_c)
    );

    fa fa_s1_c38_n78 (
        .a(stage1_col38[0]),
        .b(stage1_col38[1]),
        .c_in(stage1_col38[2]),
        .s(fa_s1_c38_n78_s),
        .c_out(fa_s1_c38_n78_c)
    );

    fa fa_s1_c38_n79 (
        .a(stage1_col38[3]),
        .b(stage1_col38[4]),
        .c_in(stage1_col38[5]),
        .s(fa_s1_c38_n79_s),
        .c_out(fa_s1_c38_n79_c)
    );

    fa fa_s1_c38_n80 (
        .a(stage1_col38[6]),
        .b(stage1_col38[7]),
        .c_in(stage1_col38[8]),
        .s(fa_s1_c38_n80_s),
        .c_out(fa_s1_c38_n80_c)
    );

    fa fa_s1_c38_n81 (
        .a(stage1_col38[9]),
        .b(stage1_col38[10]),
        .c_in(stage1_col38[11]),
        .s(fa_s1_c38_n81_s),
        .c_out(fa_s1_c38_n81_c)
    );

    fa fa_s1_c39_n82 (
        .a(stage1_col39[0]),
        .b(stage1_col39[1]),
        .c_in(stage1_col39[2]),
        .s(fa_s1_c39_n82_s),
        .c_out(fa_s1_c39_n82_c)
    );

    fa fa_s1_c39_n83 (
        .a(stage1_col39[3]),
        .b(stage1_col39[4]),
        .c_in(stage1_col39[5]),
        .s(fa_s1_c39_n83_s),
        .c_out(fa_s1_c39_n83_c)
    );

    fa fa_s1_c39_n84 (
        .a(stage1_col39[6]),
        .b(stage1_col39[7]),
        .c_in(stage1_col39[8]),
        .s(fa_s1_c39_n84_s),
        .c_out(fa_s1_c39_n84_c)
    );

    fa fa_s1_c39_n85 (
        .a(stage1_col39[9]),
        .b(stage1_col39[10]),
        .c_in(stage1_col39[11]),
        .s(fa_s1_c39_n85_s),
        .c_out(fa_s1_c39_n85_c)
    );

    fa fa_s1_c39_n86 (
        .a(stage1_col39[12]),
        .b(stage1_col39[13]),
        .c_in(stage1_col39[14]),
        .s(fa_s1_c39_n86_s),
        .c_out(fa_s1_c39_n86_c)
    );

    fa fa_s1_c40_n87 (
        .a(stage1_col40[0]),
        .b(stage1_col40[1]),
        .c_in(stage1_col40[2]),
        .s(fa_s1_c40_n87_s),
        .c_out(fa_s1_c40_n87_c)
    );

    fa fa_s1_c40_n88 (
        .a(stage1_col40[3]),
        .b(stage1_col40[4]),
        .c_in(stage1_col40[5]),
        .s(fa_s1_c40_n88_s),
        .c_out(fa_s1_c40_n88_c)
    );

    fa fa_s1_c40_n89 (
        .a(stage1_col40[6]),
        .b(stage1_col40[7]),
        .c_in(stage1_col40[8]),
        .s(fa_s1_c40_n89_s),
        .c_out(fa_s1_c40_n89_c)
    );

    fa fa_s1_c40_n90 (
        .a(stage1_col40[9]),
        .b(stage1_col40[10]),
        .c_in(stage1_col40[11]),
        .s(fa_s1_c40_n90_s),
        .c_out(fa_s1_c40_n90_c)
    );

    fa fa_s1_c41_n91 (
        .a(stage1_col41[0]),
        .b(stage1_col41[1]),
        .c_in(stage1_col41[2]),
        .s(fa_s1_c41_n91_s),
        .c_out(fa_s1_c41_n91_c)
    );

    fa fa_s1_c41_n92 (
        .a(stage1_col41[3]),
        .b(stage1_col41[4]),
        .c_in(stage1_col41[5]),
        .s(fa_s1_c41_n92_s),
        .c_out(fa_s1_c41_n92_c)
    );

    fa fa_s1_c41_n93 (
        .a(stage1_col41[6]),
        .b(stage1_col41[7]),
        .c_in(stage1_col41[8]),
        .s(fa_s1_c41_n93_s),
        .c_out(fa_s1_c41_n93_c)
    );

    fa fa_s1_c41_n94 (
        .a(stage1_col41[9]),
        .b(stage1_col41[10]),
        .c_in(stage1_col41[11]),
        .s(fa_s1_c41_n94_s),
        .c_out(fa_s1_c41_n94_c)
    );

    fa fa_s1_c42_n95 (
        .a(stage1_col42[0]),
        .b(stage1_col42[1]),
        .c_in(stage1_col42[2]),
        .s(fa_s1_c42_n95_s),
        .c_out(fa_s1_c42_n95_c)
    );

    fa fa_s1_c42_n96 (
        .a(stage1_col42[3]),
        .b(stage1_col42[4]),
        .c_in(stage1_col42[5]),
        .s(fa_s1_c42_n96_s),
        .c_out(fa_s1_c42_n96_c)
    );

    fa fa_s1_c42_n97 (
        .a(stage1_col42[6]),
        .b(stage1_col42[7]),
        .c_in(stage1_col42[8]),
        .s(fa_s1_c42_n97_s),
        .c_out(fa_s1_c42_n97_c)
    );

    fa fa_s1_c42_n98 (
        .a(stage1_col42[9]),
        .b(stage1_col42[10]),
        .c_in(stage1_col42[11]),
        .s(fa_s1_c42_n98_s),
        .c_out(fa_s1_c42_n98_c)
    );

    fa fa_s1_c42_n99 (
        .a(stage1_col42[12]),
        .b(stage1_col42[13]),
        .c_in(stage1_col42[14]),
        .s(fa_s1_c42_n99_s),
        .c_out(fa_s1_c42_n99_c)
    );

    fa fa_s1_c43_n100 (
        .a(stage1_col43[0]),
        .b(stage1_col43[1]),
        .c_in(stage1_col43[2]),
        .s(fa_s1_c43_n100_s),
        .c_out(fa_s1_c43_n100_c)
    );

    fa fa_s1_c43_n101 (
        .a(stage1_col43[3]),
        .b(stage1_col43[4]),
        .c_in(stage1_col43[5]),
        .s(fa_s1_c43_n101_s),
        .c_out(fa_s1_c43_n101_c)
    );

    fa fa_s1_c43_n102 (
        .a(stage1_col43[6]),
        .b(stage1_col43[7]),
        .c_in(stage1_col43[8]),
        .s(fa_s1_c43_n102_s),
        .c_out(fa_s1_c43_n102_c)
    );

    fa fa_s1_c43_n103 (
        .a(stage1_col43[9]),
        .b(stage1_col43[10]),
        .c_in(stage1_col43[11]),
        .s(fa_s1_c43_n103_s),
        .c_out(fa_s1_c43_n103_c)
    );

    fa fa_s1_c43_n104 (
        .a(stage1_col43[12]),
        .b(stage1_col43[13]),
        .c_in(stage1_col43[14]),
        .s(fa_s1_c43_n104_s),
        .c_out(fa_s1_c43_n104_c)
    );

    fa fa_s1_c44_n105 (
        .a(stage1_col44[0]),
        .b(stage1_col44[1]),
        .c_in(stage1_col44[2]),
        .s(fa_s1_c44_n105_s),
        .c_out(fa_s1_c44_n105_c)
    );

    fa fa_s1_c44_n106 (
        .a(stage1_col44[3]),
        .b(stage1_col44[4]),
        .c_in(stage1_col44[5]),
        .s(fa_s1_c44_n106_s),
        .c_out(fa_s1_c44_n106_c)
    );

    fa fa_s1_c44_n107 (
        .a(stage1_col44[6]),
        .b(stage1_col44[7]),
        .c_in(stage1_col44[8]),
        .s(fa_s1_c44_n107_s),
        .c_out(fa_s1_c44_n107_c)
    );

    fa fa_s1_c44_n108 (
        .a(stage1_col44[9]),
        .b(stage1_col44[10]),
        .c_in(stage1_col44[11]),
        .s(fa_s1_c44_n108_s),
        .c_out(fa_s1_c44_n108_c)
    );

    fa fa_s1_c44_n109 (
        .a(stage1_col44[12]),
        .b(stage1_col44[13]),
        .c_in(stage1_col44[14]),
        .s(fa_s1_c44_n109_s),
        .c_out(fa_s1_c44_n109_c)
    );

    fa fa_s1_c45_n110 (
        .a(stage1_col45[0]),
        .b(stage1_col45[1]),
        .c_in(stage1_col45[2]),
        .s(fa_s1_c45_n110_s),
        .c_out(fa_s1_c45_n110_c)
    );

    fa fa_s1_c45_n111 (
        .a(stage1_col45[3]),
        .b(stage1_col45[4]),
        .c_in(stage1_col45[5]),
        .s(fa_s1_c45_n111_s),
        .c_out(fa_s1_c45_n111_c)
    );

    fa fa_s1_c45_n112 (
        .a(stage1_col45[6]),
        .b(stage1_col45[7]),
        .c_in(stage1_col45[8]),
        .s(fa_s1_c45_n112_s),
        .c_out(fa_s1_c45_n112_c)
    );

    fa fa_s1_c45_n113 (
        .a(stage1_col45[9]),
        .b(stage1_col45[10]),
        .c_in(stage1_col45[11]),
        .s(fa_s1_c45_n113_s),
        .c_out(fa_s1_c45_n113_c)
    );

    fa fa_s1_c45_n114 (
        .a(stage1_col45[12]),
        .b(stage1_col45[13]),
        .c_in(stage1_col45[14]),
        .s(fa_s1_c45_n114_s),
        .c_out(fa_s1_c45_n114_c)
    );

    fa fa_s1_c46_n115 (
        .a(stage1_col46[0]),
        .b(stage1_col46[1]),
        .c_in(stage1_col46[2]),
        .s(fa_s1_c46_n115_s),
        .c_out(fa_s1_c46_n115_c)
    );

    fa fa_s1_c46_n116 (
        .a(stage1_col46[3]),
        .b(stage1_col46[4]),
        .c_in(stage1_col46[5]),
        .s(fa_s1_c46_n116_s),
        .c_out(fa_s1_c46_n116_c)
    );

    fa fa_s1_c46_n117 (
        .a(stage1_col46[6]),
        .b(stage1_col46[7]),
        .c_in(stage1_col46[8]),
        .s(fa_s1_c46_n117_s),
        .c_out(fa_s1_c46_n117_c)
    );

    fa fa_s1_c46_n118 (
        .a(stage1_col46[9]),
        .b(stage1_col46[10]),
        .c_in(stage1_col46[11]),
        .s(fa_s1_c46_n118_s),
        .c_out(fa_s1_c46_n118_c)
    );

    fa fa_s1_c46_n119 (
        .a(stage1_col46[12]),
        .b(stage1_col46[13]),
        .c_in(stage1_col46[14]),
        .s(fa_s1_c46_n119_s),
        .c_out(fa_s1_c46_n119_c)
    );

    fa fa_s1_c47_n120 (
        .a(stage1_col47[0]),
        .b(stage1_col47[1]),
        .c_in(stage1_col47[2]),
        .s(fa_s1_c47_n120_s),
        .c_out(fa_s1_c47_n120_c)
    );

    fa fa_s1_c47_n121 (
        .a(stage1_col47[3]),
        .b(stage1_col47[4]),
        .c_in(stage1_col47[5]),
        .s(fa_s1_c47_n121_s),
        .c_out(fa_s1_c47_n121_c)
    );

    fa fa_s1_c47_n122 (
        .a(stage1_col47[6]),
        .b(stage1_col47[7]),
        .c_in(stage1_col47[8]),
        .s(fa_s1_c47_n122_s),
        .c_out(fa_s1_c47_n122_c)
    );

    fa fa_s1_c47_n123 (
        .a(stage1_col47[9]),
        .b(stage1_col47[10]),
        .c_in(stage1_col47[11]),
        .s(fa_s1_c47_n123_s),
        .c_out(fa_s1_c47_n123_c)
    );

    fa fa_s1_c47_n124 (
        .a(stage1_col47[12]),
        .b(stage1_col47[13]),
        .c_in(stage1_col47[14]),
        .s(fa_s1_c47_n124_s),
        .c_out(fa_s1_c47_n124_c)
    );

    fa fa_s1_c48_n125 (
        .a(stage1_col48[0]),
        .b(stage1_col48[1]),
        .c_in(stage1_col48[2]),
        .s(fa_s1_c48_n125_s),
        .c_out(fa_s1_c48_n125_c)
    );

    fa fa_s1_c48_n126 (
        .a(stage1_col48[3]),
        .b(stage1_col48[4]),
        .c_in(stage1_col48[5]),
        .s(fa_s1_c48_n126_s),
        .c_out(fa_s1_c48_n126_c)
    );

    fa fa_s1_c48_n127 (
        .a(stage1_col48[6]),
        .b(stage1_col48[7]),
        .c_in(stage1_col48[8]),
        .s(fa_s1_c48_n127_s),
        .c_out(fa_s1_c48_n127_c)
    );

    fa fa_s1_c48_n128 (
        .a(stage1_col48[9]),
        .b(stage1_col48[10]),
        .c_in(stage1_col48[11]),
        .s(fa_s1_c48_n128_s),
        .c_out(fa_s1_c48_n128_c)
    );

    fa fa_s1_c48_n129 (
        .a(stage1_col48[12]),
        .b(stage1_col48[13]),
        .c_in(stage1_col48[14]),
        .s(fa_s1_c48_n129_s),
        .c_out(fa_s1_c48_n129_c)
    );

    fa fa_s1_c48_n130 (
        .a(stage1_col48[15]),
        .b(stage1_col48[16]),
        .c_in(stage1_col48[17]),
        .s(fa_s1_c48_n130_s),
        .c_out(fa_s1_c48_n130_c)
    );

    fa fa_s1_c49_n131 (
        .a(stage1_col49[0]),
        .b(stage1_col49[1]),
        .c_in(stage1_col49[2]),
        .s(fa_s1_c49_n131_s),
        .c_out(fa_s1_c49_n131_c)
    );

    fa fa_s1_c49_n132 (
        .a(stage1_col49[3]),
        .b(stage1_col49[4]),
        .c_in(stage1_col49[5]),
        .s(fa_s1_c49_n132_s),
        .c_out(fa_s1_c49_n132_c)
    );

    fa fa_s1_c49_n133 (
        .a(stage1_col49[6]),
        .b(stage1_col49[7]),
        .c_in(stage1_col49[8]),
        .s(fa_s1_c49_n133_s),
        .c_out(fa_s1_c49_n133_c)
    );

    fa fa_s1_c49_n134 (
        .a(stage1_col49[9]),
        .b(stage1_col49[10]),
        .c_in(stage1_col49[11]),
        .s(fa_s1_c49_n134_s),
        .c_out(fa_s1_c49_n134_c)
    );

    fa fa_s1_c49_n135 (
        .a(stage1_col49[12]),
        .b(stage1_col49[13]),
        .c_in(stage1_col49[14]),
        .s(fa_s1_c49_n135_s),
        .c_out(fa_s1_c49_n135_c)
    );

    fa fa_s1_c50_n136 (
        .a(stage1_col50[0]),
        .b(stage1_col50[1]),
        .c_in(stage1_col50[2]),
        .s(fa_s1_c50_n136_s),
        .c_out(fa_s1_c50_n136_c)
    );

    fa fa_s1_c50_n137 (
        .a(stage1_col50[3]),
        .b(stage1_col50[4]),
        .c_in(stage1_col50[5]),
        .s(fa_s1_c50_n137_s),
        .c_out(fa_s1_c50_n137_c)
    );

    fa fa_s1_c50_n138 (
        .a(stage1_col50[6]),
        .b(stage1_col50[7]),
        .c_in(stage1_col50[8]),
        .s(fa_s1_c50_n138_s),
        .c_out(fa_s1_c50_n138_c)
    );

    fa fa_s1_c50_n139 (
        .a(stage1_col50[9]),
        .b(stage1_col50[10]),
        .c_in(stage1_col50[11]),
        .s(fa_s1_c50_n139_s),
        .c_out(fa_s1_c50_n139_c)
    );

    fa fa_s1_c50_n140 (
        .a(stage1_col50[12]),
        .b(stage1_col50[13]),
        .c_in(stage1_col50[14]),
        .s(fa_s1_c50_n140_s),
        .c_out(fa_s1_c50_n140_c)
    );

    fa fa_s1_c51_n141 (
        .a(stage1_col51[0]),
        .b(stage1_col51[1]),
        .c_in(stage1_col51[2]),
        .s(fa_s1_c51_n141_s),
        .c_out(fa_s1_c51_n141_c)
    );

    fa fa_s1_c51_n142 (
        .a(stage1_col51[3]),
        .b(stage1_col51[4]),
        .c_in(stage1_col51[5]),
        .s(fa_s1_c51_n142_s),
        .c_out(fa_s1_c51_n142_c)
    );

    fa fa_s1_c51_n143 (
        .a(stage1_col51[6]),
        .b(stage1_col51[7]),
        .c_in(stage1_col51[8]),
        .s(fa_s1_c51_n143_s),
        .c_out(fa_s1_c51_n143_c)
    );

    fa fa_s1_c51_n144 (
        .a(stage1_col51[9]),
        .b(stage1_col51[10]),
        .c_in(stage1_col51[11]),
        .s(fa_s1_c51_n144_s),
        .c_out(fa_s1_c51_n144_c)
    );

    fa fa_s1_c51_n145 (
        .a(stage1_col51[12]),
        .b(stage1_col51[13]),
        .c_in(stage1_col51[14]),
        .s(fa_s1_c51_n145_s),
        .c_out(fa_s1_c51_n145_c)
    );

    fa fa_s1_c51_n146 (
        .a(stage1_col51[15]),
        .b(stage1_col51[16]),
        .c_in(stage1_col51[17]),
        .s(fa_s1_c51_n146_s),
        .c_out(fa_s1_c51_n146_c)
    );

    fa fa_s1_c52_n147 (
        .a(stage1_col52[0]),
        .b(stage1_col52[1]),
        .c_in(stage1_col52[2]),
        .s(fa_s1_c52_n147_s),
        .c_out(fa_s1_c52_n147_c)
    );

    fa fa_s1_c52_n148 (
        .a(stage1_col52[3]),
        .b(stage1_col52[4]),
        .c_in(stage1_col52[5]),
        .s(fa_s1_c52_n148_s),
        .c_out(fa_s1_c52_n148_c)
    );

    fa fa_s1_c52_n149 (
        .a(stage1_col52[6]),
        .b(stage1_col52[7]),
        .c_in(stage1_col52[8]),
        .s(fa_s1_c52_n149_s),
        .c_out(fa_s1_c52_n149_c)
    );

    fa fa_s1_c52_n150 (
        .a(stage1_col52[9]),
        .b(stage1_col52[10]),
        .c_in(stage1_col52[11]),
        .s(fa_s1_c52_n150_s),
        .c_out(fa_s1_c52_n150_c)
    );

    fa fa_s1_c52_n151 (
        .a(stage1_col52[12]),
        .b(stage1_col52[13]),
        .c_in(stage1_col52[14]),
        .s(fa_s1_c52_n151_s),
        .c_out(fa_s1_c52_n151_c)
    );

    fa fa_s1_c52_n152 (
        .a(stage1_col52[15]),
        .b(stage1_col52[16]),
        .c_in(stage1_col52[17]),
        .s(fa_s1_c52_n152_s),
        .c_out(fa_s1_c52_n152_c)
    );

    fa fa_s1_c53_n153 (
        .a(stage1_col53[0]),
        .b(stage1_col53[1]),
        .c_in(stage1_col53[2]),
        .s(fa_s1_c53_n153_s),
        .c_out(fa_s1_c53_n153_c)
    );

    fa fa_s1_c53_n154 (
        .a(stage1_col53[3]),
        .b(stage1_col53[4]),
        .c_in(stage1_col53[5]),
        .s(fa_s1_c53_n154_s),
        .c_out(fa_s1_c53_n154_c)
    );

    fa fa_s1_c53_n155 (
        .a(stage1_col53[6]),
        .b(stage1_col53[7]),
        .c_in(stage1_col53[8]),
        .s(fa_s1_c53_n155_s),
        .c_out(fa_s1_c53_n155_c)
    );

    fa fa_s1_c53_n156 (
        .a(stage1_col53[9]),
        .b(stage1_col53[10]),
        .c_in(stage1_col53[11]),
        .s(fa_s1_c53_n156_s),
        .c_out(fa_s1_c53_n156_c)
    );

    fa fa_s1_c53_n157 (
        .a(stage1_col53[12]),
        .b(stage1_col53[13]),
        .c_in(stage1_col53[14]),
        .s(fa_s1_c53_n157_s),
        .c_out(fa_s1_c53_n157_c)
    );

    fa fa_s1_c53_n158 (
        .a(stage1_col53[15]),
        .b(stage1_col53[16]),
        .c_in(stage1_col53[17]),
        .s(fa_s1_c53_n158_s),
        .c_out(fa_s1_c53_n158_c)
    );

    fa fa_s1_c54_n159 (
        .a(stage1_col54[0]),
        .b(stage1_col54[1]),
        .c_in(stage1_col54[2]),
        .s(fa_s1_c54_n159_s),
        .c_out(fa_s1_c54_n159_c)
    );

    fa fa_s1_c54_n160 (
        .a(stage1_col54[3]),
        .b(stage1_col54[4]),
        .c_in(stage1_col54[5]),
        .s(fa_s1_c54_n160_s),
        .c_out(fa_s1_c54_n160_c)
    );

    fa fa_s1_c54_n161 (
        .a(stage1_col54[6]),
        .b(stage1_col54[7]),
        .c_in(stage1_col54[8]),
        .s(fa_s1_c54_n161_s),
        .c_out(fa_s1_c54_n161_c)
    );

    fa fa_s1_c54_n162 (
        .a(stage1_col54[9]),
        .b(stage1_col54[10]),
        .c_in(stage1_col54[11]),
        .s(fa_s1_c54_n162_s),
        .c_out(fa_s1_c54_n162_c)
    );

    fa fa_s1_c54_n163 (
        .a(stage1_col54[12]),
        .b(stage1_col54[13]),
        .c_in(stage1_col54[14]),
        .s(fa_s1_c54_n163_s),
        .c_out(fa_s1_c54_n163_c)
    );

    fa fa_s1_c54_n164 (
        .a(stage1_col54[15]),
        .b(stage1_col54[16]),
        .c_in(stage1_col54[17]),
        .s(fa_s1_c54_n164_s),
        .c_out(fa_s1_c54_n164_c)
    );

    fa fa_s1_c55_n165 (
        .a(stage1_col55[0]),
        .b(stage1_col55[1]),
        .c_in(stage1_col55[2]),
        .s(fa_s1_c55_n165_s),
        .c_out(fa_s1_c55_n165_c)
    );

    fa fa_s1_c55_n166 (
        .a(stage1_col55[3]),
        .b(stage1_col55[4]),
        .c_in(stage1_col55[5]),
        .s(fa_s1_c55_n166_s),
        .c_out(fa_s1_c55_n166_c)
    );

    fa fa_s1_c55_n167 (
        .a(stage1_col55[6]),
        .b(stage1_col55[7]),
        .c_in(stage1_col55[8]),
        .s(fa_s1_c55_n167_s),
        .c_out(fa_s1_c55_n167_c)
    );

    fa fa_s1_c55_n168 (
        .a(stage1_col55[9]),
        .b(stage1_col55[10]),
        .c_in(stage1_col55[11]),
        .s(fa_s1_c55_n168_s),
        .c_out(fa_s1_c55_n168_c)
    );

    fa fa_s1_c55_n169 (
        .a(stage1_col55[12]),
        .b(stage1_col55[13]),
        .c_in(stage1_col55[14]),
        .s(fa_s1_c55_n169_s),
        .c_out(fa_s1_c55_n169_c)
    );

    fa fa_s1_c55_n170 (
        .a(stage1_col55[15]),
        .b(stage1_col55[16]),
        .c_in(stage1_col55[17]),
        .s(fa_s1_c55_n170_s),
        .c_out(fa_s1_c55_n170_c)
    );

    fa fa_s1_c56_n171 (
        .a(stage1_col56[0]),
        .b(stage1_col56[1]),
        .c_in(stage1_col56[2]),
        .s(fa_s1_c56_n171_s),
        .c_out(fa_s1_c56_n171_c)
    );

    fa fa_s1_c56_n172 (
        .a(stage1_col56[3]),
        .b(stage1_col56[4]),
        .c_in(stage1_col56[5]),
        .s(fa_s1_c56_n172_s),
        .c_out(fa_s1_c56_n172_c)
    );

    fa fa_s1_c56_n173 (
        .a(stage1_col56[6]),
        .b(stage1_col56[7]),
        .c_in(stage1_col56[8]),
        .s(fa_s1_c56_n173_s),
        .c_out(fa_s1_c56_n173_c)
    );

    fa fa_s1_c56_n174 (
        .a(stage1_col56[9]),
        .b(stage1_col56[10]),
        .c_in(stage1_col56[11]),
        .s(fa_s1_c56_n174_s),
        .c_out(fa_s1_c56_n174_c)
    );

    fa fa_s1_c56_n175 (
        .a(stage1_col56[12]),
        .b(stage1_col56[13]),
        .c_in(stage1_col56[14]),
        .s(fa_s1_c56_n175_s),
        .c_out(fa_s1_c56_n175_c)
    );

    fa fa_s1_c56_n176 (
        .a(stage1_col56[15]),
        .b(stage1_col56[16]),
        .c_in(stage1_col56[17]),
        .s(fa_s1_c56_n176_s),
        .c_out(fa_s1_c56_n176_c)
    );

    fa fa_s1_c57_n177 (
        .a(stage1_col57[0]),
        .b(stage1_col57[1]),
        .c_in(stage1_col57[2]),
        .s(fa_s1_c57_n177_s),
        .c_out(fa_s1_c57_n177_c)
    );

    fa fa_s1_c57_n178 (
        .a(stage1_col57[3]),
        .b(stage1_col57[4]),
        .c_in(stage1_col57[5]),
        .s(fa_s1_c57_n178_s),
        .c_out(fa_s1_c57_n178_c)
    );

    fa fa_s1_c57_n179 (
        .a(stage1_col57[6]),
        .b(stage1_col57[7]),
        .c_in(stage1_col57[8]),
        .s(fa_s1_c57_n179_s),
        .c_out(fa_s1_c57_n179_c)
    );

    fa fa_s1_c57_n180 (
        .a(stage1_col57[9]),
        .b(stage1_col57[10]),
        .c_in(stage1_col57[11]),
        .s(fa_s1_c57_n180_s),
        .c_out(fa_s1_c57_n180_c)
    );

    fa fa_s1_c57_n181 (
        .a(stage1_col57[12]),
        .b(stage1_col57[13]),
        .c_in(stage1_col57[14]),
        .s(fa_s1_c57_n181_s),
        .c_out(fa_s1_c57_n181_c)
    );

    fa fa_s1_c57_n182 (
        .a(stage1_col57[15]),
        .b(stage1_col57[16]),
        .c_in(stage1_col57[17]),
        .s(fa_s1_c57_n182_s),
        .c_out(fa_s1_c57_n182_c)
    );

    fa fa_s1_c57_n183 (
        .a(stage1_col57[18]),
        .b(stage1_col57[19]),
        .c_in(stage1_col57[20]),
        .s(fa_s1_c57_n183_s),
        .c_out(fa_s1_c57_n183_c)
    );

    fa fa_s1_c58_n184 (
        .a(stage1_col58[0]),
        .b(stage1_col58[1]),
        .c_in(stage1_col58[2]),
        .s(fa_s1_c58_n184_s),
        .c_out(fa_s1_c58_n184_c)
    );

    fa fa_s1_c58_n185 (
        .a(stage1_col58[3]),
        .b(stage1_col58[4]),
        .c_in(stage1_col58[5]),
        .s(fa_s1_c58_n185_s),
        .c_out(fa_s1_c58_n185_c)
    );

    fa fa_s1_c58_n186 (
        .a(stage1_col58[6]),
        .b(stage1_col58[7]),
        .c_in(stage1_col58[8]),
        .s(fa_s1_c58_n186_s),
        .c_out(fa_s1_c58_n186_c)
    );

    fa fa_s1_c58_n187 (
        .a(stage1_col58[9]),
        .b(stage1_col58[10]),
        .c_in(stage1_col58[11]),
        .s(fa_s1_c58_n187_s),
        .c_out(fa_s1_c58_n187_c)
    );

    fa fa_s1_c58_n188 (
        .a(stage1_col58[12]),
        .b(stage1_col58[13]),
        .c_in(stage1_col58[14]),
        .s(fa_s1_c58_n188_s),
        .c_out(fa_s1_c58_n188_c)
    );

    fa fa_s1_c58_n189 (
        .a(stage1_col58[15]),
        .b(stage1_col58[16]),
        .c_in(stage1_col58[17]),
        .s(fa_s1_c58_n189_s),
        .c_out(fa_s1_c58_n189_c)
    );

    fa fa_s1_c59_n190 (
        .a(stage1_col59[0]),
        .b(stage1_col59[1]),
        .c_in(stage1_col59[2]),
        .s(fa_s1_c59_n190_s),
        .c_out(fa_s1_c59_n190_c)
    );

    fa fa_s1_c59_n191 (
        .a(stage1_col59[3]),
        .b(stage1_col59[4]),
        .c_in(stage1_col59[5]),
        .s(fa_s1_c59_n191_s),
        .c_out(fa_s1_c59_n191_c)
    );

    fa fa_s1_c59_n192 (
        .a(stage1_col59[6]),
        .b(stage1_col59[7]),
        .c_in(stage1_col59[8]),
        .s(fa_s1_c59_n192_s),
        .c_out(fa_s1_c59_n192_c)
    );

    fa fa_s1_c59_n193 (
        .a(stage1_col59[9]),
        .b(stage1_col59[10]),
        .c_in(stage1_col59[11]),
        .s(fa_s1_c59_n193_s),
        .c_out(fa_s1_c59_n193_c)
    );

    fa fa_s1_c59_n194 (
        .a(stage1_col59[12]),
        .b(stage1_col59[13]),
        .c_in(stage1_col59[14]),
        .s(fa_s1_c59_n194_s),
        .c_out(fa_s1_c59_n194_c)
    );

    fa fa_s1_c59_n195 (
        .a(stage1_col59[15]),
        .b(stage1_col59[16]),
        .c_in(stage1_col59[17]),
        .s(fa_s1_c59_n195_s),
        .c_out(fa_s1_c59_n195_c)
    );

    fa fa_s1_c60_n196 (
        .a(stage1_col60[0]),
        .b(stage1_col60[1]),
        .c_in(stage1_col60[2]),
        .s(fa_s1_c60_n196_s),
        .c_out(fa_s1_c60_n196_c)
    );

    fa fa_s1_c60_n197 (
        .a(stage1_col60[3]),
        .b(stage1_col60[4]),
        .c_in(stage1_col60[5]),
        .s(fa_s1_c60_n197_s),
        .c_out(fa_s1_c60_n197_c)
    );

    fa fa_s1_c60_n198 (
        .a(stage1_col60[6]),
        .b(stage1_col60[7]),
        .c_in(stage1_col60[8]),
        .s(fa_s1_c60_n198_s),
        .c_out(fa_s1_c60_n198_c)
    );

    fa fa_s1_c60_n199 (
        .a(stage1_col60[9]),
        .b(stage1_col60[10]),
        .c_in(stage1_col60[11]),
        .s(fa_s1_c60_n199_s),
        .c_out(fa_s1_c60_n199_c)
    );

    fa fa_s1_c60_n200 (
        .a(stage1_col60[12]),
        .b(stage1_col60[13]),
        .c_in(stage1_col60[14]),
        .s(fa_s1_c60_n200_s),
        .c_out(fa_s1_c60_n200_c)
    );

    fa fa_s1_c60_n201 (
        .a(stage1_col60[15]),
        .b(stage1_col60[16]),
        .c_in(stage1_col60[17]),
        .s(fa_s1_c60_n201_s),
        .c_out(fa_s1_c60_n201_c)
    );

    fa fa_s1_c60_n202 (
        .a(stage1_col60[18]),
        .b(stage1_col60[19]),
        .c_in(stage1_col60[20]),
        .s(fa_s1_c60_n202_s),
        .c_out(fa_s1_c60_n202_c)
    );

    fa fa_s1_c61_n203 (
        .a(stage1_col61[0]),
        .b(stage1_col61[1]),
        .c_in(stage1_col61[2]),
        .s(fa_s1_c61_n203_s),
        .c_out(fa_s1_c61_n203_c)
    );

    fa fa_s1_c61_n204 (
        .a(stage1_col61[3]),
        .b(stage1_col61[4]),
        .c_in(stage1_col61[5]),
        .s(fa_s1_c61_n204_s),
        .c_out(fa_s1_c61_n204_c)
    );

    fa fa_s1_c61_n205 (
        .a(stage1_col61[6]),
        .b(stage1_col61[7]),
        .c_in(stage1_col61[8]),
        .s(fa_s1_c61_n205_s),
        .c_out(fa_s1_c61_n205_c)
    );

    fa fa_s1_c61_n206 (
        .a(stage1_col61[9]),
        .b(stage1_col61[10]),
        .c_in(stage1_col61[11]),
        .s(fa_s1_c61_n206_s),
        .c_out(fa_s1_c61_n206_c)
    );

    fa fa_s1_c61_n207 (
        .a(stage1_col61[12]),
        .b(stage1_col61[13]),
        .c_in(stage1_col61[14]),
        .s(fa_s1_c61_n207_s),
        .c_out(fa_s1_c61_n207_c)
    );

    fa fa_s1_c61_n208 (
        .a(stage1_col61[15]),
        .b(stage1_col61[16]),
        .c_in(stage1_col61[17]),
        .s(fa_s1_c61_n208_s),
        .c_out(fa_s1_c61_n208_c)
    );

    fa fa_s1_c61_n209 (
        .a(stage1_col61[18]),
        .b(stage1_col61[19]),
        .c_in(stage1_col61[20]),
        .s(fa_s1_c61_n209_s),
        .c_out(fa_s1_c61_n209_c)
    );

    fa fa_s1_c62_n210 (
        .a(stage1_col62[0]),
        .b(stage1_col62[1]),
        .c_in(stage1_col62[2]),
        .s(fa_s1_c62_n210_s),
        .c_out(fa_s1_c62_n210_c)
    );

    fa fa_s1_c62_n211 (
        .a(stage1_col62[3]),
        .b(stage1_col62[4]),
        .c_in(stage1_col62[5]),
        .s(fa_s1_c62_n211_s),
        .c_out(fa_s1_c62_n211_c)
    );

    fa fa_s1_c62_n212 (
        .a(stage1_col62[6]),
        .b(stage1_col62[7]),
        .c_in(stage1_col62[8]),
        .s(fa_s1_c62_n212_s),
        .c_out(fa_s1_c62_n212_c)
    );

    fa fa_s1_c62_n213 (
        .a(stage1_col62[9]),
        .b(stage1_col62[10]),
        .c_in(stage1_col62[11]),
        .s(fa_s1_c62_n213_s),
        .c_out(fa_s1_c62_n213_c)
    );

    fa fa_s1_c62_n214 (
        .a(stage1_col62[12]),
        .b(stage1_col62[13]),
        .c_in(stage1_col62[14]),
        .s(fa_s1_c62_n214_s),
        .c_out(fa_s1_c62_n214_c)
    );

    fa fa_s1_c62_n215 (
        .a(stage1_col62[15]),
        .b(stage1_col62[16]),
        .c_in(stage1_col62[17]),
        .s(fa_s1_c62_n215_s),
        .c_out(fa_s1_c62_n215_c)
    );

    fa fa_s1_c62_n216 (
        .a(stage1_col62[18]),
        .b(stage1_col62[19]),
        .c_in(stage1_col62[20]),
        .s(fa_s1_c62_n216_s),
        .c_out(fa_s1_c62_n216_c)
    );

    fa fa_s1_c63_n217 (
        .a(stage1_col63[0]),
        .b(stage1_col63[1]),
        .c_in(stage1_col63[2]),
        .s(fa_s1_c63_n217_s),
        .c_out(fa_s1_c63_n217_c)
    );

    fa fa_s1_c63_n218 (
        .a(stage1_col63[3]),
        .b(stage1_col63[4]),
        .c_in(stage1_col63[5]),
        .s(fa_s1_c63_n218_s),
        .c_out(fa_s1_c63_n218_c)
    );

    fa fa_s1_c63_n219 (
        .a(stage1_col63[6]),
        .b(stage1_col63[7]),
        .c_in(stage1_col63[8]),
        .s(fa_s1_c63_n219_s),
        .c_out(fa_s1_c63_n219_c)
    );

    fa fa_s1_c63_n220 (
        .a(stage1_col63[9]),
        .b(stage1_col63[10]),
        .c_in(stage1_col63[11]),
        .s(fa_s1_c63_n220_s),
        .c_out(fa_s1_c63_n220_c)
    );

    fa fa_s1_c63_n221 (
        .a(stage1_col63[12]),
        .b(stage1_col63[13]),
        .c_in(stage1_col63[14]),
        .s(fa_s1_c63_n221_s),
        .c_out(fa_s1_c63_n221_c)
    );

    fa fa_s1_c63_n222 (
        .a(stage1_col63[15]),
        .b(stage1_col63[16]),
        .c_in(stage1_col63[17]),
        .s(fa_s1_c63_n222_s),
        .c_out(fa_s1_c63_n222_c)
    );

    fa fa_s1_c63_n223 (
        .a(stage1_col63[18]),
        .b(stage1_col63[19]),
        .c_in(stage1_col63[20]),
        .s(fa_s1_c63_n223_s),
        .c_out(fa_s1_c63_n223_c)
    );

    fa fa_s1_c64_n224 (
        .a(stage1_col64[0]),
        .b(stage1_col64[1]),
        .c_in(stage1_col64[2]),
        .s(fa_s1_c64_n224_s),
        .c_out(fa_s1_c64_n224_c)
    );

    fa fa_s1_c64_n225 (
        .a(stage1_col64[3]),
        .b(stage1_col64[4]),
        .c_in(stage1_col64[5]),
        .s(fa_s1_c64_n225_s),
        .c_out(fa_s1_c64_n225_c)
    );

    fa fa_s1_c64_n226 (
        .a(stage1_col64[6]),
        .b(stage1_col64[7]),
        .c_in(stage1_col64[8]),
        .s(fa_s1_c64_n226_s),
        .c_out(fa_s1_c64_n226_c)
    );

    fa fa_s1_c64_n227 (
        .a(stage1_col64[9]),
        .b(stage1_col64[10]),
        .c_in(stage1_col64[11]),
        .s(fa_s1_c64_n227_s),
        .c_out(fa_s1_c64_n227_c)
    );

    fa fa_s1_c64_n228 (
        .a(stage1_col64[12]),
        .b(stage1_col64[13]),
        .c_in(stage1_col64[14]),
        .s(fa_s1_c64_n228_s),
        .c_out(fa_s1_c64_n228_c)
    );

    fa fa_s1_c64_n229 (
        .a(stage1_col64[15]),
        .b(stage1_col64[16]),
        .c_in(stage1_col64[17]),
        .s(fa_s1_c64_n229_s),
        .c_out(fa_s1_c64_n229_c)
    );

    fa fa_s1_c64_n230 (
        .a(stage1_col64[18]),
        .b(stage1_col64[19]),
        .c_in(stage1_col64[20]),
        .s(fa_s1_c64_n230_s),
        .c_out(fa_s1_c64_n230_c)
    );

    fa fa_s1_c65_n231 (
        .a(stage1_col65[0]),
        .b(stage1_col65[1]),
        .c_in(stage1_col65[2]),
        .s(fa_s1_c65_n231_s),
        .c_out(fa_s1_c65_n231_c)
    );

    fa fa_s1_c65_n232 (
        .a(stage1_col65[3]),
        .b(stage1_col65[4]),
        .c_in(stage1_col65[5]),
        .s(fa_s1_c65_n232_s),
        .c_out(fa_s1_c65_n232_c)
    );

    fa fa_s1_c65_n233 (
        .a(stage1_col65[6]),
        .b(stage1_col65[7]),
        .c_in(stage1_col65[8]),
        .s(fa_s1_c65_n233_s),
        .c_out(fa_s1_c65_n233_c)
    );

    fa fa_s1_c65_n234 (
        .a(stage1_col65[9]),
        .b(stage1_col65[10]),
        .c_in(stage1_col65[11]),
        .s(fa_s1_c65_n234_s),
        .c_out(fa_s1_c65_n234_c)
    );

    fa fa_s1_c65_n235 (
        .a(stage1_col65[12]),
        .b(stage1_col65[13]),
        .c_in(stage1_col65[14]),
        .s(fa_s1_c65_n235_s),
        .c_out(fa_s1_c65_n235_c)
    );

    fa fa_s1_c65_n236 (
        .a(stage1_col65[15]),
        .b(stage1_col65[16]),
        .c_in(stage1_col65[17]),
        .s(fa_s1_c65_n236_s),
        .c_out(fa_s1_c65_n236_c)
    );

    fa fa_s1_c65_n237 (
        .a(stage1_col65[18]),
        .b(stage1_col65[19]),
        .c_in(stage1_col65[20]),
        .s(fa_s1_c65_n237_s),
        .c_out(fa_s1_c65_n237_c)
    );

    fa fa_s1_c66_n238 (
        .a(stage1_col66[0]),
        .b(stage1_col66[1]),
        .c_in(stage1_col66[2]),
        .s(fa_s1_c66_n238_s),
        .c_out(fa_s1_c66_n238_c)
    );

    fa fa_s1_c66_n239 (
        .a(stage1_col66[3]),
        .b(stage1_col66[4]),
        .c_in(stage1_col66[5]),
        .s(fa_s1_c66_n239_s),
        .c_out(fa_s1_c66_n239_c)
    );

    fa fa_s1_c66_n240 (
        .a(stage1_col66[6]),
        .b(stage1_col66[7]),
        .c_in(stage1_col66[8]),
        .s(fa_s1_c66_n240_s),
        .c_out(fa_s1_c66_n240_c)
    );

    fa fa_s1_c66_n241 (
        .a(stage1_col66[9]),
        .b(stage1_col66[10]),
        .c_in(stage1_col66[11]),
        .s(fa_s1_c66_n241_s),
        .c_out(fa_s1_c66_n241_c)
    );

    fa fa_s1_c66_n242 (
        .a(stage1_col66[12]),
        .b(stage1_col66[13]),
        .c_in(stage1_col66[14]),
        .s(fa_s1_c66_n242_s),
        .c_out(fa_s1_c66_n242_c)
    );

    fa fa_s1_c66_n243 (
        .a(stage1_col66[15]),
        .b(stage1_col66[16]),
        .c_in(stage1_col66[17]),
        .s(fa_s1_c66_n243_s),
        .c_out(fa_s1_c66_n243_c)
    );

    fa fa_s1_c66_n244 (
        .a(stage1_col66[18]),
        .b(stage1_col66[19]),
        .c_in(stage1_col66[20]),
        .s(fa_s1_c66_n244_s),
        .c_out(fa_s1_c66_n244_c)
    );

    fa fa_s1_c67_n245 (
        .a(stage1_col67[0]),
        .b(stage1_col67[1]),
        .c_in(stage1_col67[2]),
        .s(fa_s1_c67_n245_s),
        .c_out(fa_s1_c67_n245_c)
    );

    fa fa_s1_c67_n246 (
        .a(stage1_col67[3]),
        .b(stage1_col67[4]),
        .c_in(stage1_col67[5]),
        .s(fa_s1_c67_n246_s),
        .c_out(fa_s1_c67_n246_c)
    );

    fa fa_s1_c67_n247 (
        .a(stage1_col67[6]),
        .b(stage1_col67[7]),
        .c_in(stage1_col67[8]),
        .s(fa_s1_c67_n247_s),
        .c_out(fa_s1_c67_n247_c)
    );

    fa fa_s1_c67_n248 (
        .a(stage1_col67[9]),
        .b(stage1_col67[10]),
        .c_in(stage1_col67[11]),
        .s(fa_s1_c67_n248_s),
        .c_out(fa_s1_c67_n248_c)
    );

    fa fa_s1_c67_n249 (
        .a(stage1_col67[12]),
        .b(stage1_col67[13]),
        .c_in(stage1_col67[14]),
        .s(fa_s1_c67_n249_s),
        .c_out(fa_s1_c67_n249_c)
    );

    fa fa_s1_c67_n250 (
        .a(stage1_col67[15]),
        .b(stage1_col67[16]),
        .c_in(stage1_col67[17]),
        .s(fa_s1_c67_n250_s),
        .c_out(fa_s1_c67_n250_c)
    );

    fa fa_s1_c67_n251 (
        .a(stage1_col67[18]),
        .b(stage1_col67[19]),
        .c_in(stage1_col67[20]),
        .s(fa_s1_c67_n251_s),
        .c_out(fa_s1_c67_n251_c)
    );

    fa fa_s1_c68_n252 (
        .a(stage1_col68[0]),
        .b(stage1_col68[1]),
        .c_in(stage1_col68[2]),
        .s(fa_s1_c68_n252_s),
        .c_out(fa_s1_c68_n252_c)
    );

    fa fa_s1_c68_n253 (
        .a(stage1_col68[3]),
        .b(stage1_col68[4]),
        .c_in(stage1_col68[5]),
        .s(fa_s1_c68_n253_s),
        .c_out(fa_s1_c68_n253_c)
    );

    fa fa_s1_c68_n254 (
        .a(stage1_col68[6]),
        .b(stage1_col68[7]),
        .c_in(stage1_col68[8]),
        .s(fa_s1_c68_n254_s),
        .c_out(fa_s1_c68_n254_c)
    );

    fa fa_s1_c68_n255 (
        .a(stage1_col68[9]),
        .b(stage1_col68[10]),
        .c_in(stage1_col68[11]),
        .s(fa_s1_c68_n255_s),
        .c_out(fa_s1_c68_n255_c)
    );

    fa fa_s1_c68_n256 (
        .a(stage1_col68[12]),
        .b(stage1_col68[13]),
        .c_in(stage1_col68[14]),
        .s(fa_s1_c68_n256_s),
        .c_out(fa_s1_c68_n256_c)
    );

    fa fa_s1_c68_n257 (
        .a(stage1_col68[15]),
        .b(stage1_col68[16]),
        .c_in(stage1_col68[17]),
        .s(fa_s1_c68_n257_s),
        .c_out(fa_s1_c68_n257_c)
    );

    fa fa_s1_c68_n258 (
        .a(stage1_col68[18]),
        .b(stage1_col68[19]),
        .c_in(stage1_col68[20]),
        .s(fa_s1_c68_n258_s),
        .c_out(fa_s1_c68_n258_c)
    );

    fa fa_s1_c69_n259 (
        .a(stage1_col69[0]),
        .b(stage1_col69[1]),
        .c_in(stage1_col69[2]),
        .s(fa_s1_c69_n259_s),
        .c_out(fa_s1_c69_n259_c)
    );

    fa fa_s1_c69_n260 (
        .a(stage1_col69[3]),
        .b(stage1_col69[4]),
        .c_in(stage1_col69[5]),
        .s(fa_s1_c69_n260_s),
        .c_out(fa_s1_c69_n260_c)
    );

    fa fa_s1_c69_n261 (
        .a(stage1_col69[6]),
        .b(stage1_col69[7]),
        .c_in(stage1_col69[8]),
        .s(fa_s1_c69_n261_s),
        .c_out(fa_s1_c69_n261_c)
    );

    fa fa_s1_c69_n262 (
        .a(stage1_col69[9]),
        .b(stage1_col69[10]),
        .c_in(stage1_col69[11]),
        .s(fa_s1_c69_n262_s),
        .c_out(fa_s1_c69_n262_c)
    );

    fa fa_s1_c69_n263 (
        .a(stage1_col69[12]),
        .b(stage1_col69[13]),
        .c_in(stage1_col69[14]),
        .s(fa_s1_c69_n263_s),
        .c_out(fa_s1_c69_n263_c)
    );

    fa fa_s1_c69_n264 (
        .a(stage1_col69[15]),
        .b(stage1_col69[16]),
        .c_in(stage1_col69[17]),
        .s(fa_s1_c69_n264_s),
        .c_out(fa_s1_c69_n264_c)
    );

    fa fa_s1_c69_n265 (
        .a(stage1_col69[18]),
        .b(stage1_col69[19]),
        .c_in(stage1_col69[20]),
        .s(fa_s1_c69_n265_s),
        .c_out(fa_s1_c69_n265_c)
    );

    fa fa_s1_c70_n266 (
        .a(stage1_col70[0]),
        .b(stage1_col70[1]),
        .c_in(stage1_col70[2]),
        .s(fa_s1_c70_n266_s),
        .c_out(fa_s1_c70_n266_c)
    );

    fa fa_s1_c70_n267 (
        .a(stage1_col70[3]),
        .b(stage1_col70[4]),
        .c_in(stage1_col70[5]),
        .s(fa_s1_c70_n267_s),
        .c_out(fa_s1_c70_n267_c)
    );

    fa fa_s1_c70_n268 (
        .a(stage1_col70[6]),
        .b(stage1_col70[7]),
        .c_in(stage1_col70[8]),
        .s(fa_s1_c70_n268_s),
        .c_out(fa_s1_c70_n268_c)
    );

    fa fa_s1_c70_n269 (
        .a(stage1_col70[9]),
        .b(stage1_col70[10]),
        .c_in(stage1_col70[11]),
        .s(fa_s1_c70_n269_s),
        .c_out(fa_s1_c70_n269_c)
    );

    fa fa_s1_c70_n270 (
        .a(stage1_col70[12]),
        .b(stage1_col70[13]),
        .c_in(stage1_col70[14]),
        .s(fa_s1_c70_n270_s),
        .c_out(fa_s1_c70_n270_c)
    );

    fa fa_s1_c70_n271 (
        .a(stage1_col70[15]),
        .b(stage1_col70[16]),
        .c_in(stage1_col70[17]),
        .s(fa_s1_c70_n271_s),
        .c_out(fa_s1_c70_n271_c)
    );

    fa fa_s1_c70_n272 (
        .a(stage1_col70[18]),
        .b(stage1_col70[19]),
        .c_in(stage1_col70[20]),
        .s(fa_s1_c70_n272_s),
        .c_out(fa_s1_c70_n272_c)
    );

    fa fa_s1_c71_n273 (
        .a(stage1_col71[0]),
        .b(stage1_col71[1]),
        .c_in(stage1_col71[2]),
        .s(fa_s1_c71_n273_s),
        .c_out(fa_s1_c71_n273_c)
    );

    fa fa_s1_c71_n274 (
        .a(stage1_col71[3]),
        .b(stage1_col71[4]),
        .c_in(stage1_col71[5]),
        .s(fa_s1_c71_n274_s),
        .c_out(fa_s1_c71_n274_c)
    );

    fa fa_s1_c71_n275 (
        .a(stage1_col71[6]),
        .b(stage1_col71[7]),
        .c_in(stage1_col71[8]),
        .s(fa_s1_c71_n275_s),
        .c_out(fa_s1_c71_n275_c)
    );

    fa fa_s1_c71_n276 (
        .a(stage1_col71[9]),
        .b(stage1_col71[10]),
        .c_in(stage1_col71[11]),
        .s(fa_s1_c71_n276_s),
        .c_out(fa_s1_c71_n276_c)
    );

    fa fa_s1_c71_n277 (
        .a(stage1_col71[12]),
        .b(stage1_col71[13]),
        .c_in(stage1_col71[14]),
        .s(fa_s1_c71_n277_s),
        .c_out(fa_s1_c71_n277_c)
    );

    fa fa_s1_c71_n278 (
        .a(stage1_col71[15]),
        .b(stage1_col71[16]),
        .c_in(stage1_col71[17]),
        .s(fa_s1_c71_n278_s),
        .c_out(fa_s1_c71_n278_c)
    );

    fa fa_s1_c71_n279 (
        .a(stage1_col71[18]),
        .b(stage1_col71[19]),
        .c_in(stage1_col71[20]),
        .s(fa_s1_c71_n279_s),
        .c_out(fa_s1_c71_n279_c)
    );

    fa fa_s1_c72_n280 (
        .a(stage1_col72[0]),
        .b(stage1_col72[1]),
        .c_in(stage1_col72[2]),
        .s(fa_s1_c72_n280_s),
        .c_out(fa_s1_c72_n280_c)
    );

    fa fa_s1_c72_n281 (
        .a(stage1_col72[3]),
        .b(stage1_col72[4]),
        .c_in(stage1_col72[5]),
        .s(fa_s1_c72_n281_s),
        .c_out(fa_s1_c72_n281_c)
    );

    fa fa_s1_c72_n282 (
        .a(stage1_col72[6]),
        .b(stage1_col72[7]),
        .c_in(stage1_col72[8]),
        .s(fa_s1_c72_n282_s),
        .c_out(fa_s1_c72_n282_c)
    );

    fa fa_s1_c72_n283 (
        .a(stage1_col72[9]),
        .b(stage1_col72[10]),
        .c_in(stage1_col72[11]),
        .s(fa_s1_c72_n283_s),
        .c_out(fa_s1_c72_n283_c)
    );

    fa fa_s1_c72_n284 (
        .a(stage1_col72[12]),
        .b(stage1_col72[13]),
        .c_in(stage1_col72[14]),
        .s(fa_s1_c72_n284_s),
        .c_out(fa_s1_c72_n284_c)
    );

    fa fa_s1_c72_n285 (
        .a(stage1_col72[15]),
        .b(stage1_col72[16]),
        .c_in(stage1_col72[17]),
        .s(fa_s1_c72_n285_s),
        .c_out(fa_s1_c72_n285_c)
    );

    fa fa_s1_c72_n286 (
        .a(stage1_col72[18]),
        .b(stage1_col72[19]),
        .c_in(stage1_col72[20]),
        .s(fa_s1_c72_n286_s),
        .c_out(fa_s1_c72_n286_c)
    );

    fa fa_s1_c73_n287 (
        .a(stage1_col73[0]),
        .b(stage1_col73[1]),
        .c_in(stage1_col73[2]),
        .s(fa_s1_c73_n287_s),
        .c_out(fa_s1_c73_n287_c)
    );

    fa fa_s1_c73_n288 (
        .a(stage1_col73[3]),
        .b(stage1_col73[4]),
        .c_in(stage1_col73[5]),
        .s(fa_s1_c73_n288_s),
        .c_out(fa_s1_c73_n288_c)
    );

    fa fa_s1_c73_n289 (
        .a(stage1_col73[6]),
        .b(stage1_col73[7]),
        .c_in(stage1_col73[8]),
        .s(fa_s1_c73_n289_s),
        .c_out(fa_s1_c73_n289_c)
    );

    fa fa_s1_c73_n290 (
        .a(stage1_col73[9]),
        .b(stage1_col73[10]),
        .c_in(stage1_col73[11]),
        .s(fa_s1_c73_n290_s),
        .c_out(fa_s1_c73_n290_c)
    );

    fa fa_s1_c73_n291 (
        .a(stage1_col73[12]),
        .b(stage1_col73[13]),
        .c_in(stage1_col73[14]),
        .s(fa_s1_c73_n291_s),
        .c_out(fa_s1_c73_n291_c)
    );

    fa fa_s1_c73_n292 (
        .a(stage1_col73[15]),
        .b(stage1_col73[16]),
        .c_in(stage1_col73[17]),
        .s(fa_s1_c73_n292_s),
        .c_out(fa_s1_c73_n292_c)
    );

    fa fa_s1_c73_n293 (
        .a(stage1_col73[18]),
        .b(stage1_col73[19]),
        .c_in(stage1_col73[20]),
        .s(fa_s1_c73_n293_s),
        .c_out(fa_s1_c73_n293_c)
    );

    fa fa_s1_c74_n294 (
        .a(stage1_col74[0]),
        .b(stage1_col74[1]),
        .c_in(stage1_col74[2]),
        .s(fa_s1_c74_n294_s),
        .c_out(fa_s1_c74_n294_c)
    );

    fa fa_s1_c74_n295 (
        .a(stage1_col74[3]),
        .b(stage1_col74[4]),
        .c_in(stage1_col74[5]),
        .s(fa_s1_c74_n295_s),
        .c_out(fa_s1_c74_n295_c)
    );

    fa fa_s1_c74_n296 (
        .a(stage1_col74[6]),
        .b(stage1_col74[7]),
        .c_in(stage1_col74[8]),
        .s(fa_s1_c74_n296_s),
        .c_out(fa_s1_c74_n296_c)
    );

    fa fa_s1_c74_n297 (
        .a(stage1_col74[9]),
        .b(stage1_col74[10]),
        .c_in(stage1_col74[11]),
        .s(fa_s1_c74_n297_s),
        .c_out(fa_s1_c74_n297_c)
    );

    fa fa_s1_c74_n298 (
        .a(stage1_col74[12]),
        .b(stage1_col74[13]),
        .c_in(stage1_col74[14]),
        .s(fa_s1_c74_n298_s),
        .c_out(fa_s1_c74_n298_c)
    );

    fa fa_s1_c74_n299 (
        .a(stage1_col74[15]),
        .b(stage1_col74[16]),
        .c_in(stage1_col74[17]),
        .s(fa_s1_c74_n299_s),
        .c_out(fa_s1_c74_n299_c)
    );

    fa fa_s1_c74_n300 (
        .a(stage1_col74[18]),
        .b(stage1_col74[19]),
        .c_in(stage1_col74[20]),
        .s(fa_s1_c74_n300_s),
        .c_out(fa_s1_c74_n300_c)
    );

    fa fa_s1_c75_n301 (
        .a(stage1_col75[0]),
        .b(stage1_col75[1]),
        .c_in(stage1_col75[2]),
        .s(fa_s1_c75_n301_s),
        .c_out(fa_s1_c75_n301_c)
    );

    fa fa_s1_c75_n302 (
        .a(stage1_col75[3]),
        .b(stage1_col75[4]),
        .c_in(stage1_col75[5]),
        .s(fa_s1_c75_n302_s),
        .c_out(fa_s1_c75_n302_c)
    );

    fa fa_s1_c75_n303 (
        .a(stage1_col75[6]),
        .b(stage1_col75[7]),
        .c_in(stage1_col75[8]),
        .s(fa_s1_c75_n303_s),
        .c_out(fa_s1_c75_n303_c)
    );

    fa fa_s1_c75_n304 (
        .a(stage1_col75[9]),
        .b(stage1_col75[10]),
        .c_in(stage1_col75[11]),
        .s(fa_s1_c75_n304_s),
        .c_out(fa_s1_c75_n304_c)
    );

    fa fa_s1_c75_n305 (
        .a(stage1_col75[12]),
        .b(stage1_col75[13]),
        .c_in(stage1_col75[14]),
        .s(fa_s1_c75_n305_s),
        .c_out(fa_s1_c75_n305_c)
    );

    fa fa_s1_c75_n306 (
        .a(stage1_col75[15]),
        .b(stage1_col75[16]),
        .c_in(stage1_col75[17]),
        .s(fa_s1_c75_n306_s),
        .c_out(fa_s1_c75_n306_c)
    );

    fa fa_s1_c75_n307 (
        .a(stage1_col75[18]),
        .b(stage1_col75[19]),
        .c_in(stage1_col75[20]),
        .s(fa_s1_c75_n307_s),
        .c_out(fa_s1_c75_n307_c)
    );

    fa fa_s1_c76_n308 (
        .a(stage1_col76[0]),
        .b(stage1_col76[1]),
        .c_in(stage1_col76[2]),
        .s(fa_s1_c76_n308_s),
        .c_out(fa_s1_c76_n308_c)
    );

    fa fa_s1_c76_n309 (
        .a(stage1_col76[3]),
        .b(stage1_col76[4]),
        .c_in(stage1_col76[5]),
        .s(fa_s1_c76_n309_s),
        .c_out(fa_s1_c76_n309_c)
    );

    fa fa_s1_c76_n310 (
        .a(stage1_col76[6]),
        .b(stage1_col76[7]),
        .c_in(stage1_col76[8]),
        .s(fa_s1_c76_n310_s),
        .c_out(fa_s1_c76_n310_c)
    );

    fa fa_s1_c76_n311 (
        .a(stage1_col76[9]),
        .b(stage1_col76[10]),
        .c_in(stage1_col76[11]),
        .s(fa_s1_c76_n311_s),
        .c_out(fa_s1_c76_n311_c)
    );

    fa fa_s1_c76_n312 (
        .a(stage1_col76[12]),
        .b(stage1_col76[13]),
        .c_in(stage1_col76[14]),
        .s(fa_s1_c76_n312_s),
        .c_out(fa_s1_c76_n312_c)
    );

    fa fa_s1_c76_n313 (
        .a(stage1_col76[15]),
        .b(stage1_col76[16]),
        .c_in(stage1_col76[17]),
        .s(fa_s1_c76_n313_s),
        .c_out(fa_s1_c76_n313_c)
    );

    fa fa_s1_c76_n314 (
        .a(stage1_col76[18]),
        .b(stage1_col76[19]),
        .c_in(stage1_col76[20]),
        .s(fa_s1_c76_n314_s),
        .c_out(fa_s1_c76_n314_c)
    );

    fa fa_s1_c77_n315 (
        .a(stage1_col77[0]),
        .b(stage1_col77[1]),
        .c_in(stage1_col77[2]),
        .s(fa_s1_c77_n315_s),
        .c_out(fa_s1_c77_n315_c)
    );

    fa fa_s1_c77_n316 (
        .a(stage1_col77[3]),
        .b(stage1_col77[4]),
        .c_in(stage1_col77[5]),
        .s(fa_s1_c77_n316_s),
        .c_out(fa_s1_c77_n316_c)
    );

    fa fa_s1_c77_n317 (
        .a(stage1_col77[6]),
        .b(stage1_col77[7]),
        .c_in(stage1_col77[8]),
        .s(fa_s1_c77_n317_s),
        .c_out(fa_s1_c77_n317_c)
    );

    fa fa_s1_c77_n318 (
        .a(stage1_col77[9]),
        .b(stage1_col77[10]),
        .c_in(stage1_col77[11]),
        .s(fa_s1_c77_n318_s),
        .c_out(fa_s1_c77_n318_c)
    );

    fa fa_s1_c77_n319 (
        .a(stage1_col77[12]),
        .b(stage1_col77[13]),
        .c_in(stage1_col77[14]),
        .s(fa_s1_c77_n319_s),
        .c_out(fa_s1_c77_n319_c)
    );

    fa fa_s1_c77_n320 (
        .a(stage1_col77[15]),
        .b(stage1_col77[16]),
        .c_in(stage1_col77[17]),
        .s(fa_s1_c77_n320_s),
        .c_out(fa_s1_c77_n320_c)
    );

    fa fa_s1_c77_n321 (
        .a(stage1_col77[18]),
        .b(stage1_col77[19]),
        .c_in(stage1_col77[20]),
        .s(fa_s1_c77_n321_s),
        .c_out(fa_s1_c77_n321_c)
    );

    fa fa_s1_c78_n322 (
        .a(stage1_col78[0]),
        .b(stage1_col78[1]),
        .c_in(stage1_col78[2]),
        .s(fa_s1_c78_n322_s),
        .c_out(fa_s1_c78_n322_c)
    );

    fa fa_s1_c78_n323 (
        .a(stage1_col78[3]),
        .b(stage1_col78[4]),
        .c_in(stage1_col78[5]),
        .s(fa_s1_c78_n323_s),
        .c_out(fa_s1_c78_n323_c)
    );

    fa fa_s1_c78_n324 (
        .a(stage1_col78[6]),
        .b(stage1_col78[7]),
        .c_in(stage1_col78[8]),
        .s(fa_s1_c78_n324_s),
        .c_out(fa_s1_c78_n324_c)
    );

    fa fa_s1_c78_n325 (
        .a(stage1_col78[9]),
        .b(stage1_col78[10]),
        .c_in(stage1_col78[11]),
        .s(fa_s1_c78_n325_s),
        .c_out(fa_s1_c78_n325_c)
    );

    fa fa_s1_c78_n326 (
        .a(stage1_col78[12]),
        .b(stage1_col78[13]),
        .c_in(stage1_col78[14]),
        .s(fa_s1_c78_n326_s),
        .c_out(fa_s1_c78_n326_c)
    );

    fa fa_s1_c78_n327 (
        .a(stage1_col78[15]),
        .b(stage1_col78[16]),
        .c_in(stage1_col78[17]),
        .s(fa_s1_c78_n327_s),
        .c_out(fa_s1_c78_n327_c)
    );

    fa fa_s1_c78_n328 (
        .a(stage1_col78[18]),
        .b(stage1_col78[19]),
        .c_in(stage1_col78[20]),
        .s(fa_s1_c78_n328_s),
        .c_out(fa_s1_c78_n328_c)
    );

    fa fa_s1_c79_n329 (
        .a(stage1_col79[0]),
        .b(stage1_col79[1]),
        .c_in(stage1_col79[2]),
        .s(fa_s1_c79_n329_s),
        .c_out(fa_s1_c79_n329_c)
    );

    fa fa_s1_c79_n330 (
        .a(stage1_col79[3]),
        .b(stage1_col79[4]),
        .c_in(stage1_col79[5]),
        .s(fa_s1_c79_n330_s),
        .c_out(fa_s1_c79_n330_c)
    );

    fa fa_s1_c79_n331 (
        .a(stage1_col79[6]),
        .b(stage1_col79[7]),
        .c_in(stage1_col79[8]),
        .s(fa_s1_c79_n331_s),
        .c_out(fa_s1_c79_n331_c)
    );

    fa fa_s1_c79_n332 (
        .a(stage1_col79[9]),
        .b(stage1_col79[10]),
        .c_in(stage1_col79[11]),
        .s(fa_s1_c79_n332_s),
        .c_out(fa_s1_c79_n332_c)
    );

    fa fa_s1_c79_n333 (
        .a(stage1_col79[12]),
        .b(stage1_col79[13]),
        .c_in(stage1_col79[14]),
        .s(fa_s1_c79_n333_s),
        .c_out(fa_s1_c79_n333_c)
    );

    fa fa_s1_c79_n334 (
        .a(stage1_col79[15]),
        .b(stage1_col79[16]),
        .c_in(stage1_col79[17]),
        .s(fa_s1_c79_n334_s),
        .c_out(fa_s1_c79_n334_c)
    );

    fa fa_s1_c79_n335 (
        .a(stage1_col79[18]),
        .b(stage1_col79[19]),
        .c_in(stage1_col79[20]),
        .s(fa_s1_c79_n335_s),
        .c_out(fa_s1_c79_n335_c)
    );

    fa fa_s1_c80_n336 (
        .a(stage1_col80[0]),
        .b(stage1_col80[1]),
        .c_in(stage1_col80[2]),
        .s(fa_s1_c80_n336_s),
        .c_out(fa_s1_c80_n336_c)
    );

    fa fa_s1_c80_n337 (
        .a(stage1_col80[3]),
        .b(stage1_col80[4]),
        .c_in(stage1_col80[5]),
        .s(fa_s1_c80_n337_s),
        .c_out(fa_s1_c80_n337_c)
    );

    fa fa_s1_c80_n338 (
        .a(stage1_col80[6]),
        .b(stage1_col80[7]),
        .c_in(stage1_col80[8]),
        .s(fa_s1_c80_n338_s),
        .c_out(fa_s1_c80_n338_c)
    );

    fa fa_s1_c80_n339 (
        .a(stage1_col80[9]),
        .b(stage1_col80[10]),
        .c_in(stage1_col80[11]),
        .s(fa_s1_c80_n339_s),
        .c_out(fa_s1_c80_n339_c)
    );

    fa fa_s1_c80_n340 (
        .a(stage1_col80[12]),
        .b(stage1_col80[13]),
        .c_in(stage1_col80[14]),
        .s(fa_s1_c80_n340_s),
        .c_out(fa_s1_c80_n340_c)
    );

    fa fa_s1_c80_n341 (
        .a(stage1_col80[15]),
        .b(stage1_col80[16]),
        .c_in(stage1_col80[17]),
        .s(fa_s1_c80_n341_s),
        .c_out(fa_s1_c80_n341_c)
    );

    fa fa_s1_c80_n342 (
        .a(stage1_col80[18]),
        .b(stage1_col80[19]),
        .c_in(stage1_col80[20]),
        .s(fa_s1_c80_n342_s),
        .c_out(fa_s1_c80_n342_c)
    );

    fa fa_s1_c81_n343 (
        .a(stage1_col81[0]),
        .b(stage1_col81[1]),
        .c_in(stage1_col81[2]),
        .s(fa_s1_c81_n343_s),
        .c_out(fa_s1_c81_n343_c)
    );

    fa fa_s1_c81_n344 (
        .a(stage1_col81[3]),
        .b(stage1_col81[4]),
        .c_in(stage1_col81[5]),
        .s(fa_s1_c81_n344_s),
        .c_out(fa_s1_c81_n344_c)
    );

    fa fa_s1_c81_n345 (
        .a(stage1_col81[6]),
        .b(stage1_col81[7]),
        .c_in(stage1_col81[8]),
        .s(fa_s1_c81_n345_s),
        .c_out(fa_s1_c81_n345_c)
    );

    fa fa_s1_c81_n346 (
        .a(stage1_col81[9]),
        .b(stage1_col81[10]),
        .c_in(stage1_col81[11]),
        .s(fa_s1_c81_n346_s),
        .c_out(fa_s1_c81_n346_c)
    );

    fa fa_s1_c81_n347 (
        .a(stage1_col81[12]),
        .b(stage1_col81[13]),
        .c_in(stage1_col81[14]),
        .s(fa_s1_c81_n347_s),
        .c_out(fa_s1_c81_n347_c)
    );

    fa fa_s1_c81_n348 (
        .a(stage1_col81[15]),
        .b(stage1_col81[16]),
        .c_in(stage1_col81[17]),
        .s(fa_s1_c81_n348_s),
        .c_out(fa_s1_c81_n348_c)
    );

    fa fa_s1_c81_n349 (
        .a(stage1_col81[18]),
        .b(stage1_col81[19]),
        .c_in(stage1_col81[20]),
        .s(fa_s1_c81_n349_s),
        .c_out(fa_s1_c81_n349_c)
    );

    fa fa_s1_c82_n350 (
        .a(stage1_col82[0]),
        .b(stage1_col82[1]),
        .c_in(stage1_col82[2]),
        .s(fa_s1_c82_n350_s),
        .c_out(fa_s1_c82_n350_c)
    );

    fa fa_s1_c82_n351 (
        .a(stage1_col82[3]),
        .b(stage1_col82[4]),
        .c_in(stage1_col82[5]),
        .s(fa_s1_c82_n351_s),
        .c_out(fa_s1_c82_n351_c)
    );

    fa fa_s1_c82_n352 (
        .a(stage1_col82[6]),
        .b(stage1_col82[7]),
        .c_in(stage1_col82[8]),
        .s(fa_s1_c82_n352_s),
        .c_out(fa_s1_c82_n352_c)
    );

    fa fa_s1_c82_n353 (
        .a(stage1_col82[9]),
        .b(stage1_col82[10]),
        .c_in(stage1_col82[11]),
        .s(fa_s1_c82_n353_s),
        .c_out(fa_s1_c82_n353_c)
    );

    fa fa_s1_c82_n354 (
        .a(stage1_col82[12]),
        .b(stage1_col82[13]),
        .c_in(stage1_col82[14]),
        .s(fa_s1_c82_n354_s),
        .c_out(fa_s1_c82_n354_c)
    );

    fa fa_s1_c82_n355 (
        .a(stage1_col82[15]),
        .b(stage1_col82[16]),
        .c_in(stage1_col82[17]),
        .s(fa_s1_c82_n355_s),
        .c_out(fa_s1_c82_n355_c)
    );

    fa fa_s1_c82_n356 (
        .a(stage1_col82[18]),
        .b(stage1_col82[19]),
        .c_in(stage1_col82[20]),
        .s(fa_s1_c82_n356_s),
        .c_out(fa_s1_c82_n356_c)
    );

    fa fa_s1_c83_n357 (
        .a(stage1_col83[0]),
        .b(stage1_col83[1]),
        .c_in(stage1_col83[2]),
        .s(fa_s1_c83_n357_s),
        .c_out(fa_s1_c83_n357_c)
    );

    fa fa_s1_c83_n358 (
        .a(stage1_col83[3]),
        .b(stage1_col83[4]),
        .c_in(stage1_col83[5]),
        .s(fa_s1_c83_n358_s),
        .c_out(fa_s1_c83_n358_c)
    );

    fa fa_s1_c83_n359 (
        .a(stage1_col83[6]),
        .b(stage1_col83[7]),
        .c_in(stage1_col83[8]),
        .s(fa_s1_c83_n359_s),
        .c_out(fa_s1_c83_n359_c)
    );

    fa fa_s1_c83_n360 (
        .a(stage1_col83[9]),
        .b(stage1_col83[10]),
        .c_in(stage1_col83[11]),
        .s(fa_s1_c83_n360_s),
        .c_out(fa_s1_c83_n360_c)
    );

    fa fa_s1_c83_n361 (
        .a(stage1_col83[12]),
        .b(stage1_col83[13]),
        .c_in(stage1_col83[14]),
        .s(fa_s1_c83_n361_s),
        .c_out(fa_s1_c83_n361_c)
    );

    fa fa_s1_c83_n362 (
        .a(stage1_col83[15]),
        .b(stage1_col83[16]),
        .c_in(stage1_col83[17]),
        .s(fa_s1_c83_n362_s),
        .c_out(fa_s1_c83_n362_c)
    );

    fa fa_s1_c83_n363 (
        .a(stage1_col83[18]),
        .b(stage1_col83[19]),
        .c_in(stage1_col83[20]),
        .s(fa_s1_c83_n363_s),
        .c_out(fa_s1_c83_n363_c)
    );

    fa fa_s1_c84_n364 (
        .a(stage1_col84[0]),
        .b(stage1_col84[1]),
        .c_in(stage1_col84[2]),
        .s(fa_s1_c84_n364_s),
        .c_out(fa_s1_c84_n364_c)
    );

    fa fa_s1_c84_n365 (
        .a(stage1_col84[3]),
        .b(stage1_col84[4]),
        .c_in(stage1_col84[5]),
        .s(fa_s1_c84_n365_s),
        .c_out(fa_s1_c84_n365_c)
    );

    fa fa_s1_c84_n366 (
        .a(stage1_col84[6]),
        .b(stage1_col84[7]),
        .c_in(stage1_col84[8]),
        .s(fa_s1_c84_n366_s),
        .c_out(fa_s1_c84_n366_c)
    );

    fa fa_s1_c84_n367 (
        .a(stage1_col84[9]),
        .b(stage1_col84[10]),
        .c_in(stage1_col84[11]),
        .s(fa_s1_c84_n367_s),
        .c_out(fa_s1_c84_n367_c)
    );

    fa fa_s1_c84_n368 (
        .a(stage1_col84[12]),
        .b(stage1_col84[13]),
        .c_in(stage1_col84[14]),
        .s(fa_s1_c84_n368_s),
        .c_out(fa_s1_c84_n368_c)
    );

    fa fa_s1_c84_n369 (
        .a(stage1_col84[15]),
        .b(stage1_col84[16]),
        .c_in(stage1_col84[17]),
        .s(fa_s1_c84_n369_s),
        .c_out(fa_s1_c84_n369_c)
    );

    fa fa_s1_c84_n370 (
        .a(stage1_col84[18]),
        .b(stage1_col84[19]),
        .c_in(stage1_col84[20]),
        .s(fa_s1_c84_n370_s),
        .c_out(fa_s1_c84_n370_c)
    );

    fa fa_s1_c85_n371 (
        .a(stage1_col85[0]),
        .b(stage1_col85[1]),
        .c_in(stage1_col85[2]),
        .s(fa_s1_c85_n371_s),
        .c_out(fa_s1_c85_n371_c)
    );

    fa fa_s1_c85_n372 (
        .a(stage1_col85[3]),
        .b(stage1_col85[4]),
        .c_in(stage1_col85[5]),
        .s(fa_s1_c85_n372_s),
        .c_out(fa_s1_c85_n372_c)
    );

    fa fa_s1_c85_n373 (
        .a(stage1_col85[6]),
        .b(stage1_col85[7]),
        .c_in(stage1_col85[8]),
        .s(fa_s1_c85_n373_s),
        .c_out(fa_s1_c85_n373_c)
    );

    fa fa_s1_c85_n374 (
        .a(stage1_col85[9]),
        .b(stage1_col85[10]),
        .c_in(stage1_col85[11]),
        .s(fa_s1_c85_n374_s),
        .c_out(fa_s1_c85_n374_c)
    );

    fa fa_s1_c85_n375 (
        .a(stage1_col85[12]),
        .b(stage1_col85[13]),
        .c_in(stage1_col85[14]),
        .s(fa_s1_c85_n375_s),
        .c_out(fa_s1_c85_n375_c)
    );

    fa fa_s1_c85_n376 (
        .a(stage1_col85[15]),
        .b(stage1_col85[16]),
        .c_in(stage1_col85[17]),
        .s(fa_s1_c85_n376_s),
        .c_out(fa_s1_c85_n376_c)
    );

    fa fa_s1_c85_n377 (
        .a(stage1_col85[18]),
        .b(stage1_col85[19]),
        .c_in(stage1_col85[20]),
        .s(fa_s1_c85_n377_s),
        .c_out(fa_s1_c85_n377_c)
    );

    fa fa_s1_c86_n378 (
        .a(stage1_col86[0]),
        .b(stage1_col86[1]),
        .c_in(stage1_col86[2]),
        .s(fa_s1_c86_n378_s),
        .c_out(fa_s1_c86_n378_c)
    );

    fa fa_s1_c86_n379 (
        .a(stage1_col86[3]),
        .b(stage1_col86[4]),
        .c_in(stage1_col86[5]),
        .s(fa_s1_c86_n379_s),
        .c_out(fa_s1_c86_n379_c)
    );

    fa fa_s1_c86_n380 (
        .a(stage1_col86[6]),
        .b(stage1_col86[7]),
        .c_in(stage1_col86[8]),
        .s(fa_s1_c86_n380_s),
        .c_out(fa_s1_c86_n380_c)
    );

    fa fa_s1_c86_n381 (
        .a(stage1_col86[9]),
        .b(stage1_col86[10]),
        .c_in(stage1_col86[11]),
        .s(fa_s1_c86_n381_s),
        .c_out(fa_s1_c86_n381_c)
    );

    fa fa_s1_c86_n382 (
        .a(stage1_col86[12]),
        .b(stage1_col86[13]),
        .c_in(stage1_col86[14]),
        .s(fa_s1_c86_n382_s),
        .c_out(fa_s1_c86_n382_c)
    );

    fa fa_s1_c86_n383 (
        .a(stage1_col86[15]),
        .b(stage1_col86[16]),
        .c_in(stage1_col86[17]),
        .s(fa_s1_c86_n383_s),
        .c_out(fa_s1_c86_n383_c)
    );

    fa fa_s1_c86_n384 (
        .a(stage1_col86[18]),
        .b(stage1_col86[19]),
        .c_in(stage1_col86[20]),
        .s(fa_s1_c86_n384_s),
        .c_out(fa_s1_c86_n384_c)
    );

    fa fa_s1_c87_n385 (
        .a(stage1_col87[0]),
        .b(stage1_col87[1]),
        .c_in(stage1_col87[2]),
        .s(fa_s1_c87_n385_s),
        .c_out(fa_s1_c87_n385_c)
    );

    fa fa_s1_c87_n386 (
        .a(stage1_col87[3]),
        .b(stage1_col87[4]),
        .c_in(stage1_col87[5]),
        .s(fa_s1_c87_n386_s),
        .c_out(fa_s1_c87_n386_c)
    );

    fa fa_s1_c87_n387 (
        .a(stage1_col87[6]),
        .b(stage1_col87[7]),
        .c_in(stage1_col87[8]),
        .s(fa_s1_c87_n387_s),
        .c_out(fa_s1_c87_n387_c)
    );

    fa fa_s1_c87_n388 (
        .a(stage1_col87[9]),
        .b(stage1_col87[10]),
        .c_in(stage1_col87[11]),
        .s(fa_s1_c87_n388_s),
        .c_out(fa_s1_c87_n388_c)
    );

    fa fa_s1_c87_n389 (
        .a(stage1_col87[12]),
        .b(stage1_col87[13]),
        .c_in(stage1_col87[14]),
        .s(fa_s1_c87_n389_s),
        .c_out(fa_s1_c87_n389_c)
    );

    fa fa_s1_c87_n390 (
        .a(stage1_col87[15]),
        .b(stage1_col87[16]),
        .c_in(stage1_col87[17]),
        .s(fa_s1_c87_n390_s),
        .c_out(fa_s1_c87_n390_c)
    );

    fa fa_s1_c87_n391 (
        .a(stage1_col87[18]),
        .b(stage1_col87[19]),
        .c_in(stage1_col87[20]),
        .s(fa_s1_c87_n391_s),
        .c_out(fa_s1_c87_n391_c)
    );

    fa fa_s1_c88_n392 (
        .a(stage1_col88[0]),
        .b(stage1_col88[1]),
        .c_in(stage1_col88[2]),
        .s(fa_s1_c88_n392_s),
        .c_out(fa_s1_c88_n392_c)
    );

    fa fa_s1_c88_n393 (
        .a(stage1_col88[3]),
        .b(stage1_col88[4]),
        .c_in(stage1_col88[5]),
        .s(fa_s1_c88_n393_s),
        .c_out(fa_s1_c88_n393_c)
    );

    fa fa_s1_c88_n394 (
        .a(stage1_col88[6]),
        .b(stage1_col88[7]),
        .c_in(stage1_col88[8]),
        .s(fa_s1_c88_n394_s),
        .c_out(fa_s1_c88_n394_c)
    );

    fa fa_s1_c88_n395 (
        .a(stage1_col88[9]),
        .b(stage1_col88[10]),
        .c_in(stage1_col88[11]),
        .s(fa_s1_c88_n395_s),
        .c_out(fa_s1_c88_n395_c)
    );

    fa fa_s1_c88_n396 (
        .a(stage1_col88[12]),
        .b(stage1_col88[13]),
        .c_in(stage1_col88[14]),
        .s(fa_s1_c88_n396_s),
        .c_out(fa_s1_c88_n396_c)
    );

    fa fa_s1_c88_n397 (
        .a(stage1_col88[15]),
        .b(stage1_col88[16]),
        .c_in(stage1_col88[17]),
        .s(fa_s1_c88_n397_s),
        .c_out(fa_s1_c88_n397_c)
    );

    fa fa_s1_c88_n398 (
        .a(stage1_col88[18]),
        .b(stage1_col88[19]),
        .c_in(stage1_col88[20]),
        .s(fa_s1_c88_n398_s),
        .c_out(fa_s1_c88_n398_c)
    );

    fa fa_s1_c89_n399 (
        .a(stage1_col89[0]),
        .b(stage1_col89[1]),
        .c_in(stage1_col89[2]),
        .s(fa_s1_c89_n399_s),
        .c_out(fa_s1_c89_n399_c)
    );

    fa fa_s1_c89_n400 (
        .a(stage1_col89[3]),
        .b(stage1_col89[4]),
        .c_in(stage1_col89[5]),
        .s(fa_s1_c89_n400_s),
        .c_out(fa_s1_c89_n400_c)
    );

    fa fa_s1_c89_n401 (
        .a(stage1_col89[6]),
        .b(stage1_col89[7]),
        .c_in(stage1_col89[8]),
        .s(fa_s1_c89_n401_s),
        .c_out(fa_s1_c89_n401_c)
    );

    fa fa_s1_c89_n402 (
        .a(stage1_col89[9]),
        .b(stage1_col89[10]),
        .c_in(stage1_col89[11]),
        .s(fa_s1_c89_n402_s),
        .c_out(fa_s1_c89_n402_c)
    );

    fa fa_s1_c89_n403 (
        .a(stage1_col89[12]),
        .b(stage1_col89[13]),
        .c_in(stage1_col89[14]),
        .s(fa_s1_c89_n403_s),
        .c_out(fa_s1_c89_n403_c)
    );

    fa fa_s1_c89_n404 (
        .a(stage1_col89[15]),
        .b(stage1_col89[16]),
        .c_in(stage1_col89[17]),
        .s(fa_s1_c89_n404_s),
        .c_out(fa_s1_c89_n404_c)
    );

    fa fa_s1_c89_n405 (
        .a(stage1_col89[18]),
        .b(stage1_col89[19]),
        .c_in(stage1_col89[20]),
        .s(fa_s1_c89_n405_s),
        .c_out(fa_s1_c89_n405_c)
    );

    fa fa_s1_c90_n406 (
        .a(stage1_col90[0]),
        .b(stage1_col90[1]),
        .c_in(stage1_col90[2]),
        .s(fa_s1_c90_n406_s),
        .c_out(fa_s1_c90_n406_c)
    );

    fa fa_s1_c90_n407 (
        .a(stage1_col90[3]),
        .b(stage1_col90[4]),
        .c_in(stage1_col90[5]),
        .s(fa_s1_c90_n407_s),
        .c_out(fa_s1_c90_n407_c)
    );

    fa fa_s1_c90_n408 (
        .a(stage1_col90[6]),
        .b(stage1_col90[7]),
        .c_in(stage1_col90[8]),
        .s(fa_s1_c90_n408_s),
        .c_out(fa_s1_c90_n408_c)
    );

    fa fa_s1_c90_n409 (
        .a(stage1_col90[9]),
        .b(stage1_col90[10]),
        .c_in(stage1_col90[11]),
        .s(fa_s1_c90_n409_s),
        .c_out(fa_s1_c90_n409_c)
    );

    fa fa_s1_c90_n410 (
        .a(stage1_col90[12]),
        .b(stage1_col90[13]),
        .c_in(stage1_col90[14]),
        .s(fa_s1_c90_n410_s),
        .c_out(fa_s1_c90_n410_c)
    );

    fa fa_s1_c90_n411 (
        .a(stage1_col90[15]),
        .b(stage1_col90[16]),
        .c_in(stage1_col90[17]),
        .s(fa_s1_c90_n411_s),
        .c_out(fa_s1_c90_n411_c)
    );

    fa fa_s1_c90_n412 (
        .a(stage1_col90[18]),
        .b(stage1_col90[19]),
        .c_in(stage1_col90[20]),
        .s(fa_s1_c90_n412_s),
        .c_out(fa_s1_c90_n412_c)
    );

    fa fa_s1_c91_n413 (
        .a(stage1_col91[0]),
        .b(stage1_col91[1]),
        .c_in(stage1_col91[2]),
        .s(fa_s1_c91_n413_s),
        .c_out(fa_s1_c91_n413_c)
    );

    fa fa_s1_c91_n414 (
        .a(stage1_col91[3]),
        .b(stage1_col91[4]),
        .c_in(stage1_col91[5]),
        .s(fa_s1_c91_n414_s),
        .c_out(fa_s1_c91_n414_c)
    );

    fa fa_s1_c91_n415 (
        .a(stage1_col91[6]),
        .b(stage1_col91[7]),
        .c_in(stage1_col91[8]),
        .s(fa_s1_c91_n415_s),
        .c_out(fa_s1_c91_n415_c)
    );

    fa fa_s1_c91_n416 (
        .a(stage1_col91[9]),
        .b(stage1_col91[10]),
        .c_in(stage1_col91[11]),
        .s(fa_s1_c91_n416_s),
        .c_out(fa_s1_c91_n416_c)
    );

    fa fa_s1_c91_n417 (
        .a(stage1_col91[12]),
        .b(stage1_col91[13]),
        .c_in(stage1_col91[14]),
        .s(fa_s1_c91_n417_s),
        .c_out(fa_s1_c91_n417_c)
    );

    fa fa_s1_c91_n418 (
        .a(stage1_col91[15]),
        .b(stage1_col91[16]),
        .c_in(stage1_col91[17]),
        .s(fa_s1_c91_n418_s),
        .c_out(fa_s1_c91_n418_c)
    );

    fa fa_s1_c91_n419 (
        .a(stage1_col91[18]),
        .b(stage1_col91[19]),
        .c_in(stage1_col91[20]),
        .s(fa_s1_c91_n419_s),
        .c_out(fa_s1_c91_n419_c)
    );

    fa fa_s1_c92_n420 (
        .a(stage1_col92[0]),
        .b(stage1_col92[1]),
        .c_in(stage1_col92[2]),
        .s(fa_s1_c92_n420_s),
        .c_out(fa_s1_c92_n420_c)
    );

    fa fa_s1_c92_n421 (
        .a(stage1_col92[3]),
        .b(stage1_col92[4]),
        .c_in(stage1_col92[5]),
        .s(fa_s1_c92_n421_s),
        .c_out(fa_s1_c92_n421_c)
    );

    fa fa_s1_c92_n422 (
        .a(stage1_col92[6]),
        .b(stage1_col92[7]),
        .c_in(stage1_col92[8]),
        .s(fa_s1_c92_n422_s),
        .c_out(fa_s1_c92_n422_c)
    );

    fa fa_s1_c92_n423 (
        .a(stage1_col92[9]),
        .b(stage1_col92[10]),
        .c_in(stage1_col92[11]),
        .s(fa_s1_c92_n423_s),
        .c_out(fa_s1_c92_n423_c)
    );

    fa fa_s1_c92_n424 (
        .a(stage1_col92[12]),
        .b(stage1_col92[13]),
        .c_in(stage1_col92[14]),
        .s(fa_s1_c92_n424_s),
        .c_out(fa_s1_c92_n424_c)
    );

    fa fa_s1_c92_n425 (
        .a(stage1_col92[15]),
        .b(stage1_col92[16]),
        .c_in(stage1_col92[17]),
        .s(fa_s1_c92_n425_s),
        .c_out(fa_s1_c92_n425_c)
    );

    fa fa_s1_c92_n426 (
        .a(stage1_col92[18]),
        .b(stage1_col92[19]),
        .c_in(stage1_col92[20]),
        .s(fa_s1_c92_n426_s),
        .c_out(fa_s1_c92_n426_c)
    );

    fa fa_s1_c93_n427 (
        .a(stage1_col93[0]),
        .b(stage1_col93[1]),
        .c_in(stage1_col93[2]),
        .s(fa_s1_c93_n427_s),
        .c_out(fa_s1_c93_n427_c)
    );

    fa fa_s1_c93_n428 (
        .a(stage1_col93[3]),
        .b(stage1_col93[4]),
        .c_in(stage1_col93[5]),
        .s(fa_s1_c93_n428_s),
        .c_out(fa_s1_c93_n428_c)
    );

    fa fa_s1_c93_n429 (
        .a(stage1_col93[6]),
        .b(stage1_col93[7]),
        .c_in(stage1_col93[8]),
        .s(fa_s1_c93_n429_s),
        .c_out(fa_s1_c93_n429_c)
    );

    fa fa_s1_c93_n430 (
        .a(stage1_col93[9]),
        .b(stage1_col93[10]),
        .c_in(stage1_col93[11]),
        .s(fa_s1_c93_n430_s),
        .c_out(fa_s1_c93_n430_c)
    );

    fa fa_s1_c93_n431 (
        .a(stage1_col93[12]),
        .b(stage1_col93[13]),
        .c_in(stage1_col93[14]),
        .s(fa_s1_c93_n431_s),
        .c_out(fa_s1_c93_n431_c)
    );

    fa fa_s1_c93_n432 (
        .a(stage1_col93[15]),
        .b(stage1_col93[16]),
        .c_in(stage1_col93[17]),
        .s(fa_s1_c93_n432_s),
        .c_out(fa_s1_c93_n432_c)
    );

    fa fa_s1_c93_n433 (
        .a(stage1_col93[18]),
        .b(stage1_col93[19]),
        .c_in(stage1_col93[20]),
        .s(fa_s1_c93_n433_s),
        .c_out(fa_s1_c93_n433_c)
    );

    fa fa_s1_c94_n434 (
        .a(stage1_col94[0]),
        .b(stage1_col94[1]),
        .c_in(stage1_col94[2]),
        .s(fa_s1_c94_n434_s),
        .c_out(fa_s1_c94_n434_c)
    );

    fa fa_s1_c94_n435 (
        .a(stage1_col94[3]),
        .b(stage1_col94[4]),
        .c_in(stage1_col94[5]),
        .s(fa_s1_c94_n435_s),
        .c_out(fa_s1_c94_n435_c)
    );

    fa fa_s1_c94_n436 (
        .a(stage1_col94[6]),
        .b(stage1_col94[7]),
        .c_in(stage1_col94[8]),
        .s(fa_s1_c94_n436_s),
        .c_out(fa_s1_c94_n436_c)
    );

    fa fa_s1_c94_n437 (
        .a(stage1_col94[9]),
        .b(stage1_col94[10]),
        .c_in(stage1_col94[11]),
        .s(fa_s1_c94_n437_s),
        .c_out(fa_s1_c94_n437_c)
    );

    fa fa_s1_c94_n438 (
        .a(stage1_col94[12]),
        .b(stage1_col94[13]),
        .c_in(stage1_col94[14]),
        .s(fa_s1_c94_n438_s),
        .c_out(fa_s1_c94_n438_c)
    );

    fa fa_s1_c94_n439 (
        .a(stage1_col94[15]),
        .b(stage1_col94[16]),
        .c_in(stage1_col94[17]),
        .s(fa_s1_c94_n439_s),
        .c_out(fa_s1_c94_n439_c)
    );

    fa fa_s1_c94_n440 (
        .a(stage1_col94[18]),
        .b(stage1_col94[19]),
        .c_in(stage1_col94[20]),
        .s(fa_s1_c94_n440_s),
        .c_out(fa_s1_c94_n440_c)
    );

    fa fa_s1_c95_n441 (
        .a(stage1_col95[0]),
        .b(stage1_col95[1]),
        .c_in(stage1_col95[2]),
        .s(fa_s1_c95_n441_s),
        .c_out(fa_s1_c95_n441_c)
    );

    fa fa_s1_c95_n442 (
        .a(stage1_col95[3]),
        .b(stage1_col95[4]),
        .c_in(stage1_col95[5]),
        .s(fa_s1_c95_n442_s),
        .c_out(fa_s1_c95_n442_c)
    );

    fa fa_s1_c95_n443 (
        .a(stage1_col95[6]),
        .b(stage1_col95[7]),
        .c_in(stage1_col95[8]),
        .s(fa_s1_c95_n443_s),
        .c_out(fa_s1_c95_n443_c)
    );

    fa fa_s1_c95_n444 (
        .a(stage1_col95[9]),
        .b(stage1_col95[10]),
        .c_in(stage1_col95[11]),
        .s(fa_s1_c95_n444_s),
        .c_out(fa_s1_c95_n444_c)
    );

    fa fa_s1_c95_n445 (
        .a(stage1_col95[12]),
        .b(stage1_col95[13]),
        .c_in(stage1_col95[14]),
        .s(fa_s1_c95_n445_s),
        .c_out(fa_s1_c95_n445_c)
    );

    fa fa_s1_c95_n446 (
        .a(stage1_col95[15]),
        .b(stage1_col95[16]),
        .c_in(stage1_col95[17]),
        .s(fa_s1_c95_n446_s),
        .c_out(fa_s1_c95_n446_c)
    );

    fa fa_s1_c95_n447 (
        .a(stage1_col95[18]),
        .b(stage1_col95[19]),
        .c_in(stage1_col95[20]),
        .s(fa_s1_c95_n447_s),
        .c_out(fa_s1_c95_n447_c)
    );

    fa fa_s1_c96_n448 (
        .a(stage1_col96[0]),
        .b(stage1_col96[1]),
        .c_in(stage1_col96[2]),
        .s(fa_s1_c96_n448_s),
        .c_out(fa_s1_c96_n448_c)
    );

    fa fa_s1_c96_n449 (
        .a(stage1_col96[3]),
        .b(stage1_col96[4]),
        .c_in(stage1_col96[5]),
        .s(fa_s1_c96_n449_s),
        .c_out(fa_s1_c96_n449_c)
    );

    fa fa_s1_c96_n450 (
        .a(stage1_col96[6]),
        .b(stage1_col96[7]),
        .c_in(stage1_col96[8]),
        .s(fa_s1_c96_n450_s),
        .c_out(fa_s1_c96_n450_c)
    );

    fa fa_s1_c96_n451 (
        .a(stage1_col96[9]),
        .b(stage1_col96[10]),
        .c_in(stage1_col96[11]),
        .s(fa_s1_c96_n451_s),
        .c_out(fa_s1_c96_n451_c)
    );

    fa fa_s1_c96_n452 (
        .a(stage1_col96[12]),
        .b(stage1_col96[13]),
        .c_in(stage1_col96[14]),
        .s(fa_s1_c96_n452_s),
        .c_out(fa_s1_c96_n452_c)
    );

    fa fa_s1_c96_n453 (
        .a(stage1_col96[15]),
        .b(stage1_col96[16]),
        .c_in(stage1_col96[17]),
        .s(fa_s1_c96_n453_s),
        .c_out(fa_s1_c96_n453_c)
    );

    fa fa_s1_c96_n454 (
        .a(stage1_col96[18]),
        .b(stage1_col96[19]),
        .c_in(stage1_col96[20]),
        .s(fa_s1_c96_n454_s),
        .c_out(fa_s1_c96_n454_c)
    );

    fa fa_s1_c97_n455 (
        .a(stage1_col97[0]),
        .b(stage1_col97[1]),
        .c_in(stage1_col97[2]),
        .s(fa_s1_c97_n455_s),
        .c_out(fa_s1_c97_n455_c)
    );

    fa fa_s1_c97_n456 (
        .a(stage1_col97[3]),
        .b(stage1_col97[4]),
        .c_in(stage1_col97[5]),
        .s(fa_s1_c97_n456_s),
        .c_out(fa_s1_c97_n456_c)
    );

    fa fa_s1_c97_n457 (
        .a(stage1_col97[6]),
        .b(stage1_col97[7]),
        .c_in(stage1_col97[8]),
        .s(fa_s1_c97_n457_s),
        .c_out(fa_s1_c97_n457_c)
    );

    fa fa_s1_c97_n458 (
        .a(stage1_col97[9]),
        .b(stage1_col97[10]),
        .c_in(stage1_col97[11]),
        .s(fa_s1_c97_n458_s),
        .c_out(fa_s1_c97_n458_c)
    );

    fa fa_s1_c97_n459 (
        .a(stage1_col97[12]),
        .b(stage1_col97[13]),
        .c_in(stage1_col97[14]),
        .s(fa_s1_c97_n459_s),
        .c_out(fa_s1_c97_n459_c)
    );

    fa fa_s1_c97_n460 (
        .a(stage1_col97[15]),
        .b(stage1_col97[16]),
        .c_in(stage1_col97[17]),
        .s(fa_s1_c97_n460_s),
        .c_out(fa_s1_c97_n460_c)
    );

    fa fa_s1_c97_n461 (
        .a(stage1_col97[18]),
        .b(stage1_col97[19]),
        .c_in(stage1_col97[20]),
        .s(fa_s1_c97_n461_s),
        .c_out(fa_s1_c97_n461_c)
    );

    fa fa_s1_c98_n462 (
        .a(stage1_col98[0]),
        .b(stage1_col98[1]),
        .c_in(stage1_col98[2]),
        .s(fa_s1_c98_n462_s),
        .c_out(fa_s1_c98_n462_c)
    );

    fa fa_s1_c98_n463 (
        .a(stage1_col98[3]),
        .b(stage1_col98[4]),
        .c_in(stage1_col98[5]),
        .s(fa_s1_c98_n463_s),
        .c_out(fa_s1_c98_n463_c)
    );

    fa fa_s1_c98_n464 (
        .a(stage1_col98[6]),
        .b(stage1_col98[7]),
        .c_in(stage1_col98[8]),
        .s(fa_s1_c98_n464_s),
        .c_out(fa_s1_c98_n464_c)
    );

    fa fa_s1_c98_n465 (
        .a(stage1_col98[9]),
        .b(stage1_col98[10]),
        .c_in(stage1_col98[11]),
        .s(fa_s1_c98_n465_s),
        .c_out(fa_s1_c98_n465_c)
    );

    fa fa_s1_c98_n466 (
        .a(stage1_col98[12]),
        .b(stage1_col98[13]),
        .c_in(stage1_col98[14]),
        .s(fa_s1_c98_n466_s),
        .c_out(fa_s1_c98_n466_c)
    );

    fa fa_s1_c98_n467 (
        .a(stage1_col98[15]),
        .b(stage1_col98[16]),
        .c_in(stage1_col98[17]),
        .s(fa_s1_c98_n467_s),
        .c_out(fa_s1_c98_n467_c)
    );

    fa fa_s1_c98_n468 (
        .a(stage1_col98[18]),
        .b(stage1_col98[19]),
        .c_in(stage1_col98[20]),
        .s(fa_s1_c98_n468_s),
        .c_out(fa_s1_c98_n468_c)
    );

    fa fa_s1_c99_n469 (
        .a(stage1_col99[0]),
        .b(stage1_col99[1]),
        .c_in(stage1_col99[2]),
        .s(fa_s1_c99_n469_s),
        .c_out(fa_s1_c99_n469_c)
    );

    fa fa_s1_c99_n470 (
        .a(stage1_col99[3]),
        .b(stage1_col99[4]),
        .c_in(stage1_col99[5]),
        .s(fa_s1_c99_n470_s),
        .c_out(fa_s1_c99_n470_c)
    );

    fa fa_s1_c99_n471 (
        .a(stage1_col99[6]),
        .b(stage1_col99[7]),
        .c_in(stage1_col99[8]),
        .s(fa_s1_c99_n471_s),
        .c_out(fa_s1_c99_n471_c)
    );

    fa fa_s1_c99_n472 (
        .a(stage1_col99[9]),
        .b(stage1_col99[10]),
        .c_in(stage1_col99[11]),
        .s(fa_s1_c99_n472_s),
        .c_out(fa_s1_c99_n472_c)
    );

    fa fa_s1_c99_n473 (
        .a(stage1_col99[12]),
        .b(stage1_col99[13]),
        .c_in(stage1_col99[14]),
        .s(fa_s1_c99_n473_s),
        .c_out(fa_s1_c99_n473_c)
    );

    fa fa_s1_c99_n474 (
        .a(stage1_col99[15]),
        .b(stage1_col99[16]),
        .c_in(stage1_col99[17]),
        .s(fa_s1_c99_n474_s),
        .c_out(fa_s1_c99_n474_c)
    );

    fa fa_s1_c99_n475 (
        .a(stage1_col99[18]),
        .b(stage1_col99[19]),
        .c_in(stage1_col99[20]),
        .s(fa_s1_c99_n475_s),
        .c_out(fa_s1_c99_n475_c)
    );

    fa fa_s1_c100_n476 (
        .a(stage1_col100[0]),
        .b(stage1_col100[1]),
        .c_in(stage1_col100[2]),
        .s(fa_s1_c100_n476_s),
        .c_out(fa_s1_c100_n476_c)
    );

    fa fa_s1_c100_n477 (
        .a(stage1_col100[3]),
        .b(stage1_col100[4]),
        .c_in(stage1_col100[5]),
        .s(fa_s1_c100_n477_s),
        .c_out(fa_s1_c100_n477_c)
    );

    fa fa_s1_c100_n478 (
        .a(stage1_col100[6]),
        .b(stage1_col100[7]),
        .c_in(stage1_col100[8]),
        .s(fa_s1_c100_n478_s),
        .c_out(fa_s1_c100_n478_c)
    );

    fa fa_s1_c100_n479 (
        .a(stage1_col100[9]),
        .b(stage1_col100[10]),
        .c_in(stage1_col100[11]),
        .s(fa_s1_c100_n479_s),
        .c_out(fa_s1_c100_n479_c)
    );

    fa fa_s1_c100_n480 (
        .a(stage1_col100[12]),
        .b(stage1_col100[13]),
        .c_in(stage1_col100[14]),
        .s(fa_s1_c100_n480_s),
        .c_out(fa_s1_c100_n480_c)
    );

    fa fa_s1_c100_n481 (
        .a(stage1_col100[15]),
        .b(stage1_col100[16]),
        .c_in(stage1_col100[17]),
        .s(fa_s1_c100_n481_s),
        .c_out(fa_s1_c100_n481_c)
    );

    fa fa_s1_c100_n482 (
        .a(stage1_col100[18]),
        .b(stage1_col100[19]),
        .c_in(stage1_col100[20]),
        .s(fa_s1_c100_n482_s),
        .c_out(fa_s1_c100_n482_c)
    );

    fa fa_s1_c101_n483 (
        .a(stage1_col101[0]),
        .b(stage1_col101[1]),
        .c_in(stage1_col101[2]),
        .s(fa_s1_c101_n483_s),
        .c_out(fa_s1_c101_n483_c)
    );

    fa fa_s1_c101_n484 (
        .a(stage1_col101[3]),
        .b(stage1_col101[4]),
        .c_in(stage1_col101[5]),
        .s(fa_s1_c101_n484_s),
        .c_out(fa_s1_c101_n484_c)
    );

    fa fa_s1_c101_n485 (
        .a(stage1_col101[6]),
        .b(stage1_col101[7]),
        .c_in(stage1_col101[8]),
        .s(fa_s1_c101_n485_s),
        .c_out(fa_s1_c101_n485_c)
    );

    fa fa_s1_c101_n486 (
        .a(stage1_col101[9]),
        .b(stage1_col101[10]),
        .c_in(stage1_col101[11]),
        .s(fa_s1_c101_n486_s),
        .c_out(fa_s1_c101_n486_c)
    );

    fa fa_s1_c101_n487 (
        .a(stage1_col101[12]),
        .b(stage1_col101[13]),
        .c_in(stage1_col101[14]),
        .s(fa_s1_c101_n487_s),
        .c_out(fa_s1_c101_n487_c)
    );

    fa fa_s1_c101_n488 (
        .a(stage1_col101[15]),
        .b(stage1_col101[16]),
        .c_in(stage1_col101[17]),
        .s(fa_s1_c101_n488_s),
        .c_out(fa_s1_c101_n488_c)
    );

    fa fa_s1_c101_n489 (
        .a(stage1_col101[18]),
        .b(stage1_col101[19]),
        .c_in(stage1_col101[20]),
        .s(fa_s1_c101_n489_s),
        .c_out(fa_s1_c101_n489_c)
    );

    fa fa_s1_c102_n490 (
        .a(stage1_col102[0]),
        .b(stage1_col102[1]),
        .c_in(stage1_col102[2]),
        .s(fa_s1_c102_n490_s),
        .c_out(fa_s1_c102_n490_c)
    );

    fa fa_s1_c102_n491 (
        .a(stage1_col102[3]),
        .b(stage1_col102[4]),
        .c_in(stage1_col102[5]),
        .s(fa_s1_c102_n491_s),
        .c_out(fa_s1_c102_n491_c)
    );

    fa fa_s1_c102_n492 (
        .a(stage1_col102[6]),
        .b(stage1_col102[7]),
        .c_in(stage1_col102[8]),
        .s(fa_s1_c102_n492_s),
        .c_out(fa_s1_c102_n492_c)
    );

    fa fa_s1_c102_n493 (
        .a(stage1_col102[9]),
        .b(stage1_col102[10]),
        .c_in(stage1_col102[11]),
        .s(fa_s1_c102_n493_s),
        .c_out(fa_s1_c102_n493_c)
    );

    fa fa_s1_c102_n494 (
        .a(stage1_col102[12]),
        .b(stage1_col102[13]),
        .c_in(stage1_col102[14]),
        .s(fa_s1_c102_n494_s),
        .c_out(fa_s1_c102_n494_c)
    );

    fa fa_s1_c102_n495 (
        .a(stage1_col102[15]),
        .b(stage1_col102[16]),
        .c_in(stage1_col102[17]),
        .s(fa_s1_c102_n495_s),
        .c_out(fa_s1_c102_n495_c)
    );

    fa fa_s1_c102_n496 (
        .a(stage1_col102[18]),
        .b(stage1_col102[19]),
        .c_in(stage1_col102[20]),
        .s(fa_s1_c102_n496_s),
        .c_out(fa_s1_c102_n496_c)
    );

    fa fa_s1_c103_n497 (
        .a(stage1_col103[0]),
        .b(stage1_col103[1]),
        .c_in(stage1_col103[2]),
        .s(fa_s1_c103_n497_s),
        .c_out(fa_s1_c103_n497_c)
    );

    fa fa_s1_c103_n498 (
        .a(stage1_col103[3]),
        .b(stage1_col103[4]),
        .c_in(stage1_col103[5]),
        .s(fa_s1_c103_n498_s),
        .c_out(fa_s1_c103_n498_c)
    );

    fa fa_s1_c103_n499 (
        .a(stage1_col103[6]),
        .b(stage1_col103[7]),
        .c_in(stage1_col103[8]),
        .s(fa_s1_c103_n499_s),
        .c_out(fa_s1_c103_n499_c)
    );

    fa fa_s1_c103_n500 (
        .a(stage1_col103[9]),
        .b(stage1_col103[10]),
        .c_in(stage1_col103[11]),
        .s(fa_s1_c103_n500_s),
        .c_out(fa_s1_c103_n500_c)
    );

    fa fa_s1_c103_n501 (
        .a(stage1_col103[12]),
        .b(stage1_col103[13]),
        .c_in(stage1_col103[14]),
        .s(fa_s1_c103_n501_s),
        .c_out(fa_s1_c103_n501_c)
    );

    fa fa_s1_c103_n502 (
        .a(stage1_col103[15]),
        .b(stage1_col103[16]),
        .c_in(stage1_col103[17]),
        .s(fa_s1_c103_n502_s),
        .c_out(fa_s1_c103_n502_c)
    );

    fa fa_s1_c103_n503 (
        .a(stage1_col103[18]),
        .b(stage1_col103[19]),
        .c_in(stage1_col103[20]),
        .s(fa_s1_c103_n503_s),
        .c_out(fa_s1_c103_n503_c)
    );

    fa fa_s1_c104_n504 (
        .a(stage1_col104[0]),
        .b(stage1_col104[1]),
        .c_in(stage1_col104[2]),
        .s(fa_s1_c104_n504_s),
        .c_out(fa_s1_c104_n504_c)
    );

    fa fa_s1_c104_n505 (
        .a(stage1_col104[3]),
        .b(stage1_col104[4]),
        .c_in(stage1_col104[5]),
        .s(fa_s1_c104_n505_s),
        .c_out(fa_s1_c104_n505_c)
    );

    fa fa_s1_c104_n506 (
        .a(stage1_col104[6]),
        .b(stage1_col104[7]),
        .c_in(stage1_col104[8]),
        .s(fa_s1_c104_n506_s),
        .c_out(fa_s1_c104_n506_c)
    );

    fa fa_s1_c104_n507 (
        .a(stage1_col104[9]),
        .b(stage1_col104[10]),
        .c_in(stage1_col104[11]),
        .s(fa_s1_c104_n507_s),
        .c_out(fa_s1_c104_n507_c)
    );

    fa fa_s1_c104_n508 (
        .a(stage1_col104[12]),
        .b(stage1_col104[13]),
        .c_in(stage1_col104[14]),
        .s(fa_s1_c104_n508_s),
        .c_out(fa_s1_c104_n508_c)
    );

    fa fa_s1_c104_n509 (
        .a(stage1_col104[15]),
        .b(stage1_col104[16]),
        .c_in(stage1_col104[17]),
        .s(fa_s1_c104_n509_s),
        .c_out(fa_s1_c104_n509_c)
    );

    fa fa_s1_c104_n510 (
        .a(stage1_col104[18]),
        .b(stage1_col104[19]),
        .c_in(stage1_col104[20]),
        .s(fa_s1_c104_n510_s),
        .c_out(fa_s1_c104_n510_c)
    );

    fa fa_s1_c105_n511 (
        .a(stage1_col105[0]),
        .b(stage1_col105[1]),
        .c_in(stage1_col105[2]),
        .s(fa_s1_c105_n511_s),
        .c_out(fa_s1_c105_n511_c)
    );

    fa fa_s1_c105_n512 (
        .a(stage1_col105[3]),
        .b(stage1_col105[4]),
        .c_in(stage1_col105[5]),
        .s(fa_s1_c105_n512_s),
        .c_out(fa_s1_c105_n512_c)
    );

    fa fa_s1_c105_n513 (
        .a(stage1_col105[6]),
        .b(stage1_col105[7]),
        .c_in(stage1_col105[8]),
        .s(fa_s1_c105_n513_s),
        .c_out(fa_s1_c105_n513_c)
    );

    fa fa_s1_c105_n514 (
        .a(stage1_col105[9]),
        .b(stage1_col105[10]),
        .c_in(stage1_col105[11]),
        .s(fa_s1_c105_n514_s),
        .c_out(fa_s1_c105_n514_c)
    );

    fa fa_s1_c105_n515 (
        .a(stage1_col105[12]),
        .b(stage1_col105[13]),
        .c_in(stage1_col105[14]),
        .s(fa_s1_c105_n515_s),
        .c_out(fa_s1_c105_n515_c)
    );

    fa fa_s1_c105_n516 (
        .a(stage1_col105[15]),
        .b(stage1_col105[16]),
        .c_in(stage1_col105[17]),
        .s(fa_s1_c105_n516_s),
        .c_out(fa_s1_c105_n516_c)
    );

    fa fa_s1_c105_n517 (
        .a(stage1_col105[18]),
        .b(stage1_col105[19]),
        .c_in(stage1_col105[20]),
        .s(fa_s1_c105_n517_s),
        .c_out(fa_s1_c105_n517_c)
    );

    fa fa_s1_c106_n518 (
        .a(stage1_col106[0]),
        .b(stage1_col106[1]),
        .c_in(stage1_col106[2]),
        .s(fa_s1_c106_n518_s),
        .c_out(fa_s1_c106_n518_c)
    );

    fa fa_s1_c106_n519 (
        .a(stage1_col106[3]),
        .b(stage1_col106[4]),
        .c_in(stage1_col106[5]),
        .s(fa_s1_c106_n519_s),
        .c_out(fa_s1_c106_n519_c)
    );

    fa fa_s1_c106_n520 (
        .a(stage1_col106[6]),
        .b(stage1_col106[7]),
        .c_in(stage1_col106[8]),
        .s(fa_s1_c106_n520_s),
        .c_out(fa_s1_c106_n520_c)
    );

    fa fa_s1_c106_n521 (
        .a(stage1_col106[9]),
        .b(stage1_col106[10]),
        .c_in(stage1_col106[11]),
        .s(fa_s1_c106_n521_s),
        .c_out(fa_s1_c106_n521_c)
    );

    fa fa_s1_c106_n522 (
        .a(stage1_col106[12]),
        .b(stage1_col106[13]),
        .c_in(stage1_col106[14]),
        .s(fa_s1_c106_n522_s),
        .c_out(fa_s1_c106_n522_c)
    );

    fa fa_s1_c106_n523 (
        .a(stage1_col106[15]),
        .b(stage1_col106[16]),
        .c_in(stage1_col106[17]),
        .s(fa_s1_c106_n523_s),
        .c_out(fa_s1_c106_n523_c)
    );

    fa fa_s1_c106_n524 (
        .a(stage1_col106[18]),
        .b(stage1_col106[19]),
        .c_in(stage1_col106[20]),
        .s(fa_s1_c106_n524_s),
        .c_out(fa_s1_c106_n524_c)
    );

    fa fa_s1_c107_n525 (
        .a(stage1_col107[0]),
        .b(stage1_col107[1]),
        .c_in(stage1_col107[2]),
        .s(fa_s1_c107_n525_s),
        .c_out(fa_s1_c107_n525_c)
    );

    fa fa_s1_c107_n526 (
        .a(stage1_col107[3]),
        .b(stage1_col107[4]),
        .c_in(stage1_col107[5]),
        .s(fa_s1_c107_n526_s),
        .c_out(fa_s1_c107_n526_c)
    );

    fa fa_s1_c107_n527 (
        .a(stage1_col107[6]),
        .b(stage1_col107[7]),
        .c_in(stage1_col107[8]),
        .s(fa_s1_c107_n527_s),
        .c_out(fa_s1_c107_n527_c)
    );

    fa fa_s1_c107_n528 (
        .a(stage1_col107[9]),
        .b(stage1_col107[10]),
        .c_in(stage1_col107[11]),
        .s(fa_s1_c107_n528_s),
        .c_out(fa_s1_c107_n528_c)
    );

    fa fa_s1_c107_n529 (
        .a(stage1_col107[12]),
        .b(stage1_col107[13]),
        .c_in(stage1_col107[14]),
        .s(fa_s1_c107_n529_s),
        .c_out(fa_s1_c107_n529_c)
    );

    fa fa_s1_c107_n530 (
        .a(stage1_col107[15]),
        .b(stage1_col107[16]),
        .c_in(stage1_col107[17]),
        .s(fa_s1_c107_n530_s),
        .c_out(fa_s1_c107_n530_c)
    );

    fa fa_s1_c107_n531 (
        .a(stage1_col107[18]),
        .b(stage1_col107[19]),
        .c_in(stage1_col107[20]),
        .s(fa_s1_c107_n531_s),
        .c_out(fa_s1_c107_n531_c)
    );

    fa fa_s1_c108_n532 (
        .a(stage1_col108[0]),
        .b(stage1_col108[1]),
        .c_in(stage1_col108[2]),
        .s(fa_s1_c108_n532_s),
        .c_out(fa_s1_c108_n532_c)
    );

    fa fa_s1_c108_n533 (
        .a(stage1_col108[3]),
        .b(stage1_col108[4]),
        .c_in(stage1_col108[5]),
        .s(fa_s1_c108_n533_s),
        .c_out(fa_s1_c108_n533_c)
    );

    fa fa_s1_c108_n534 (
        .a(stage1_col108[6]),
        .b(stage1_col108[7]),
        .c_in(stage1_col108[8]),
        .s(fa_s1_c108_n534_s),
        .c_out(fa_s1_c108_n534_c)
    );

    fa fa_s1_c108_n535 (
        .a(stage1_col108[9]),
        .b(stage1_col108[10]),
        .c_in(stage1_col108[11]),
        .s(fa_s1_c108_n535_s),
        .c_out(fa_s1_c108_n535_c)
    );

    fa fa_s1_c108_n536 (
        .a(stage1_col108[12]),
        .b(stage1_col108[13]),
        .c_in(stage1_col108[14]),
        .s(fa_s1_c108_n536_s),
        .c_out(fa_s1_c108_n536_c)
    );

    fa fa_s1_c108_n537 (
        .a(stage1_col108[15]),
        .b(stage1_col108[16]),
        .c_in(stage1_col108[17]),
        .s(fa_s1_c108_n537_s),
        .c_out(fa_s1_c108_n537_c)
    );

    fa fa_s1_c108_n538 (
        .a(stage1_col108[18]),
        .b(stage1_col108[19]),
        .c_in(stage1_col108[20]),
        .s(fa_s1_c108_n538_s),
        .c_out(fa_s1_c108_n538_c)
    );

    fa fa_s1_c109_n539 (
        .a(stage1_col109[0]),
        .b(stage1_col109[1]),
        .c_in(stage1_col109[2]),
        .s(fa_s1_c109_n539_s),
        .c_out(fa_s1_c109_n539_c)
    );

    fa fa_s1_c109_n540 (
        .a(stage1_col109[3]),
        .b(stage1_col109[4]),
        .c_in(stage1_col109[5]),
        .s(fa_s1_c109_n540_s),
        .c_out(fa_s1_c109_n540_c)
    );

    fa fa_s1_c109_n541 (
        .a(stage1_col109[6]),
        .b(stage1_col109[7]),
        .c_in(stage1_col109[8]),
        .s(fa_s1_c109_n541_s),
        .c_out(fa_s1_c109_n541_c)
    );

    fa fa_s1_c109_n542 (
        .a(stage1_col109[9]),
        .b(stage1_col109[10]),
        .c_in(stage1_col109[11]),
        .s(fa_s1_c109_n542_s),
        .c_out(fa_s1_c109_n542_c)
    );

    fa fa_s1_c109_n543 (
        .a(stage1_col109[12]),
        .b(stage1_col109[13]),
        .c_in(stage1_col109[14]),
        .s(fa_s1_c109_n543_s),
        .c_out(fa_s1_c109_n543_c)
    );

    fa fa_s1_c109_n544 (
        .a(stage1_col109[15]),
        .b(stage1_col109[16]),
        .c_in(stage1_col109[17]),
        .s(fa_s1_c109_n544_s),
        .c_out(fa_s1_c109_n544_c)
    );

    fa fa_s1_c109_n545 (
        .a(stage1_col109[18]),
        .b(stage1_col109[19]),
        .c_in(stage1_col109[20]),
        .s(fa_s1_c109_n545_s),
        .c_out(fa_s1_c109_n545_c)
    );

    fa fa_s1_c110_n546 (
        .a(stage1_col110[0]),
        .b(stage1_col110[1]),
        .c_in(stage1_col110[2]),
        .s(fa_s1_c110_n546_s),
        .c_out(fa_s1_c110_n546_c)
    );

    fa fa_s1_c110_n547 (
        .a(stage1_col110[3]),
        .b(stage1_col110[4]),
        .c_in(stage1_col110[5]),
        .s(fa_s1_c110_n547_s),
        .c_out(fa_s1_c110_n547_c)
    );

    fa fa_s1_c110_n548 (
        .a(stage1_col110[6]),
        .b(stage1_col110[7]),
        .c_in(stage1_col110[8]),
        .s(fa_s1_c110_n548_s),
        .c_out(fa_s1_c110_n548_c)
    );

    fa fa_s1_c110_n549 (
        .a(stage1_col110[9]),
        .b(stage1_col110[10]),
        .c_in(stage1_col110[11]),
        .s(fa_s1_c110_n549_s),
        .c_out(fa_s1_c110_n549_c)
    );

    fa fa_s1_c110_n550 (
        .a(stage1_col110[12]),
        .b(stage1_col110[13]),
        .c_in(stage1_col110[14]),
        .s(fa_s1_c110_n550_s),
        .c_out(fa_s1_c110_n550_c)
    );

    fa fa_s1_c110_n551 (
        .a(stage1_col110[15]),
        .b(stage1_col110[16]),
        .c_in(stage1_col110[17]),
        .s(fa_s1_c110_n551_s),
        .c_out(fa_s1_c110_n551_c)
    );

    fa fa_s1_c110_n552 (
        .a(stage1_col110[18]),
        .b(stage1_col110[19]),
        .c_in(stage1_col110[20]),
        .s(fa_s1_c110_n552_s),
        .c_out(fa_s1_c110_n552_c)
    );

    fa fa_s1_c111_n553 (
        .a(stage1_col111[0]),
        .b(stage1_col111[1]),
        .c_in(stage1_col111[2]),
        .s(fa_s1_c111_n553_s),
        .c_out(fa_s1_c111_n553_c)
    );

    fa fa_s1_c111_n554 (
        .a(stage1_col111[3]),
        .b(stage1_col111[4]),
        .c_in(stage1_col111[5]),
        .s(fa_s1_c111_n554_s),
        .c_out(fa_s1_c111_n554_c)
    );

    fa fa_s1_c111_n555 (
        .a(stage1_col111[6]),
        .b(stage1_col111[7]),
        .c_in(stage1_col111[8]),
        .s(fa_s1_c111_n555_s),
        .c_out(fa_s1_c111_n555_c)
    );

    fa fa_s1_c111_n556 (
        .a(stage1_col111[9]),
        .b(stage1_col111[10]),
        .c_in(stage1_col111[11]),
        .s(fa_s1_c111_n556_s),
        .c_out(fa_s1_c111_n556_c)
    );

    fa fa_s1_c111_n557 (
        .a(stage1_col111[12]),
        .b(stage1_col111[13]),
        .c_in(stage1_col111[14]),
        .s(fa_s1_c111_n557_s),
        .c_out(fa_s1_c111_n557_c)
    );

    fa fa_s1_c111_n558 (
        .a(stage1_col111[15]),
        .b(stage1_col111[16]),
        .c_in(stage1_col111[17]),
        .s(fa_s1_c111_n558_s),
        .c_out(fa_s1_c111_n558_c)
    );

    fa fa_s1_c111_n559 (
        .a(stage1_col111[18]),
        .b(stage1_col111[19]),
        .c_in(stage1_col111[20]),
        .s(fa_s1_c111_n559_s),
        .c_out(fa_s1_c111_n559_c)
    );

    fa fa_s1_c112_n560 (
        .a(stage1_col112[0]),
        .b(stage1_col112[1]),
        .c_in(stage1_col112[2]),
        .s(fa_s1_c112_n560_s),
        .c_out(fa_s1_c112_n560_c)
    );

    fa fa_s1_c112_n561 (
        .a(stage1_col112[3]),
        .b(stage1_col112[4]),
        .c_in(stage1_col112[5]),
        .s(fa_s1_c112_n561_s),
        .c_out(fa_s1_c112_n561_c)
    );

    fa fa_s1_c112_n562 (
        .a(stage1_col112[6]),
        .b(stage1_col112[7]),
        .c_in(stage1_col112[8]),
        .s(fa_s1_c112_n562_s),
        .c_out(fa_s1_c112_n562_c)
    );

    fa fa_s1_c112_n563 (
        .a(stage1_col112[9]),
        .b(stage1_col112[10]),
        .c_in(stage1_col112[11]),
        .s(fa_s1_c112_n563_s),
        .c_out(fa_s1_c112_n563_c)
    );

    fa fa_s1_c112_n564 (
        .a(stage1_col112[12]),
        .b(stage1_col112[13]),
        .c_in(stage1_col112[14]),
        .s(fa_s1_c112_n564_s),
        .c_out(fa_s1_c112_n564_c)
    );

    fa fa_s1_c112_n565 (
        .a(stage1_col112[15]),
        .b(stage1_col112[16]),
        .c_in(stage1_col112[17]),
        .s(fa_s1_c112_n565_s),
        .c_out(fa_s1_c112_n565_c)
    );

    fa fa_s1_c112_n566 (
        .a(stage1_col112[18]),
        .b(stage1_col112[19]),
        .c_in(stage1_col112[20]),
        .s(fa_s1_c112_n566_s),
        .c_out(fa_s1_c112_n566_c)
    );

    fa fa_s1_c113_n567 (
        .a(stage1_col113[0]),
        .b(stage1_col113[1]),
        .c_in(stage1_col113[2]),
        .s(fa_s1_c113_n567_s),
        .c_out(fa_s1_c113_n567_c)
    );

    fa fa_s1_c113_n568 (
        .a(stage1_col113[3]),
        .b(stage1_col113[4]),
        .c_in(stage1_col113[5]),
        .s(fa_s1_c113_n568_s),
        .c_out(fa_s1_c113_n568_c)
    );

    fa fa_s1_c113_n569 (
        .a(stage1_col113[6]),
        .b(stage1_col113[7]),
        .c_in(stage1_col113[8]),
        .s(fa_s1_c113_n569_s),
        .c_out(fa_s1_c113_n569_c)
    );

    fa fa_s1_c113_n570 (
        .a(stage1_col113[9]),
        .b(stage1_col113[10]),
        .c_in(stage1_col113[11]),
        .s(fa_s1_c113_n570_s),
        .c_out(fa_s1_c113_n570_c)
    );

    fa fa_s1_c113_n571 (
        .a(stage1_col113[12]),
        .b(stage1_col113[13]),
        .c_in(stage1_col113[14]),
        .s(fa_s1_c113_n571_s),
        .c_out(fa_s1_c113_n571_c)
    );

    fa fa_s1_c113_n572 (
        .a(stage1_col113[15]),
        .b(stage1_col113[16]),
        .c_in(stage1_col113[17]),
        .s(fa_s1_c113_n572_s),
        .c_out(fa_s1_c113_n572_c)
    );

    fa fa_s1_c113_n573 (
        .a(stage1_col113[18]),
        .b(stage1_col113[19]),
        .c_in(stage1_col113[20]),
        .s(fa_s1_c113_n573_s),
        .c_out(fa_s1_c113_n573_c)
    );

    fa fa_s1_c114_n574 (
        .a(stage1_col114[0]),
        .b(stage1_col114[1]),
        .c_in(stage1_col114[2]),
        .s(fa_s1_c114_n574_s),
        .c_out(fa_s1_c114_n574_c)
    );

    fa fa_s1_c114_n575 (
        .a(stage1_col114[3]),
        .b(stage1_col114[4]),
        .c_in(stage1_col114[5]),
        .s(fa_s1_c114_n575_s),
        .c_out(fa_s1_c114_n575_c)
    );

    fa fa_s1_c114_n576 (
        .a(stage1_col114[6]),
        .b(stage1_col114[7]),
        .c_in(stage1_col114[8]),
        .s(fa_s1_c114_n576_s),
        .c_out(fa_s1_c114_n576_c)
    );

    fa fa_s1_c114_n577 (
        .a(stage1_col114[9]),
        .b(stage1_col114[10]),
        .c_in(stage1_col114[11]),
        .s(fa_s1_c114_n577_s),
        .c_out(fa_s1_c114_n577_c)
    );

    fa fa_s1_c114_n578 (
        .a(stage1_col114[12]),
        .b(stage1_col114[13]),
        .c_in(stage1_col114[14]),
        .s(fa_s1_c114_n578_s),
        .c_out(fa_s1_c114_n578_c)
    );

    fa fa_s1_c114_n579 (
        .a(stage1_col114[15]),
        .b(stage1_col114[16]),
        .c_in(stage1_col114[17]),
        .s(fa_s1_c114_n579_s),
        .c_out(fa_s1_c114_n579_c)
    );

    fa fa_s1_c114_n580 (
        .a(stage1_col114[18]),
        .b(stage1_col114[19]),
        .c_in(stage1_col114[20]),
        .s(fa_s1_c114_n580_s),
        .c_out(fa_s1_c114_n580_c)
    );

    fa fa_s1_c115_n581 (
        .a(stage1_col115[0]),
        .b(stage1_col115[1]),
        .c_in(stage1_col115[2]),
        .s(fa_s1_c115_n581_s),
        .c_out(fa_s1_c115_n581_c)
    );

    fa fa_s1_c115_n582 (
        .a(stage1_col115[3]),
        .b(stage1_col115[4]),
        .c_in(stage1_col115[5]),
        .s(fa_s1_c115_n582_s),
        .c_out(fa_s1_c115_n582_c)
    );

    fa fa_s1_c115_n583 (
        .a(stage1_col115[6]),
        .b(stage1_col115[7]),
        .c_in(stage1_col115[8]),
        .s(fa_s1_c115_n583_s),
        .c_out(fa_s1_c115_n583_c)
    );

    fa fa_s1_c115_n584 (
        .a(stage1_col115[9]),
        .b(stage1_col115[10]),
        .c_in(stage1_col115[11]),
        .s(fa_s1_c115_n584_s),
        .c_out(fa_s1_c115_n584_c)
    );

    fa fa_s1_c115_n585 (
        .a(stage1_col115[12]),
        .b(stage1_col115[13]),
        .c_in(stage1_col115[14]),
        .s(fa_s1_c115_n585_s),
        .c_out(fa_s1_c115_n585_c)
    );

    fa fa_s1_c115_n586 (
        .a(stage1_col115[15]),
        .b(stage1_col115[16]),
        .c_in(stage1_col115[17]),
        .s(fa_s1_c115_n586_s),
        .c_out(fa_s1_c115_n586_c)
    );

    fa fa_s1_c115_n587 (
        .a(stage1_col115[18]),
        .b(stage1_col115[19]),
        .c_in(stage1_col115[20]),
        .s(fa_s1_c115_n587_s),
        .c_out(fa_s1_c115_n587_c)
    );

    fa fa_s1_c116_n588 (
        .a(stage1_col116[0]),
        .b(stage1_col116[1]),
        .c_in(stage1_col116[2]),
        .s(fa_s1_c116_n588_s),
        .c_out(fa_s1_c116_n588_c)
    );

    fa fa_s1_c116_n589 (
        .a(stage1_col116[3]),
        .b(stage1_col116[4]),
        .c_in(stage1_col116[5]),
        .s(fa_s1_c116_n589_s),
        .c_out(fa_s1_c116_n589_c)
    );

    fa fa_s1_c116_n590 (
        .a(stage1_col116[6]),
        .b(stage1_col116[7]),
        .c_in(stage1_col116[8]),
        .s(fa_s1_c116_n590_s),
        .c_out(fa_s1_c116_n590_c)
    );

    fa fa_s1_c116_n591 (
        .a(stage1_col116[9]),
        .b(stage1_col116[10]),
        .c_in(stage1_col116[11]),
        .s(fa_s1_c116_n591_s),
        .c_out(fa_s1_c116_n591_c)
    );

    fa fa_s1_c116_n592 (
        .a(stage1_col116[12]),
        .b(stage1_col116[13]),
        .c_in(stage1_col116[14]),
        .s(fa_s1_c116_n592_s),
        .c_out(fa_s1_c116_n592_c)
    );

    fa fa_s1_c116_n593 (
        .a(stage1_col116[15]),
        .b(stage1_col116[16]),
        .c_in(stage1_col116[17]),
        .s(fa_s1_c116_n593_s),
        .c_out(fa_s1_c116_n593_c)
    );

    fa fa_s1_c116_n594 (
        .a(stage1_col116[18]),
        .b(stage1_col116[19]),
        .c_in(stage1_col116[20]),
        .s(fa_s1_c116_n594_s),
        .c_out(fa_s1_c116_n594_c)
    );

    fa fa_s1_c117_n595 (
        .a(stage1_col117[0]),
        .b(stage1_col117[1]),
        .c_in(stage1_col117[2]),
        .s(fa_s1_c117_n595_s),
        .c_out(fa_s1_c117_n595_c)
    );

    fa fa_s1_c117_n596 (
        .a(stage1_col117[3]),
        .b(stage1_col117[4]),
        .c_in(stage1_col117[5]),
        .s(fa_s1_c117_n596_s),
        .c_out(fa_s1_c117_n596_c)
    );

    fa fa_s1_c117_n597 (
        .a(stage1_col117[6]),
        .b(stage1_col117[7]),
        .c_in(stage1_col117[8]),
        .s(fa_s1_c117_n597_s),
        .c_out(fa_s1_c117_n597_c)
    );

    fa fa_s1_c117_n598 (
        .a(stage1_col117[9]),
        .b(stage1_col117[10]),
        .c_in(stage1_col117[11]),
        .s(fa_s1_c117_n598_s),
        .c_out(fa_s1_c117_n598_c)
    );

    fa fa_s1_c117_n599 (
        .a(stage1_col117[12]),
        .b(stage1_col117[13]),
        .c_in(stage1_col117[14]),
        .s(fa_s1_c117_n599_s),
        .c_out(fa_s1_c117_n599_c)
    );

    fa fa_s1_c117_n600 (
        .a(stage1_col117[15]),
        .b(stage1_col117[16]),
        .c_in(stage1_col117[17]),
        .s(fa_s1_c117_n600_s),
        .c_out(fa_s1_c117_n600_c)
    );

    fa fa_s1_c117_n601 (
        .a(stage1_col117[18]),
        .b(stage1_col117[19]),
        .c_in(stage1_col117[20]),
        .s(fa_s1_c117_n601_s),
        .c_out(fa_s1_c117_n601_c)
    );

    fa fa_s1_c118_n602 (
        .a(stage1_col118[0]),
        .b(stage1_col118[1]),
        .c_in(stage1_col118[2]),
        .s(fa_s1_c118_n602_s),
        .c_out(fa_s1_c118_n602_c)
    );

    fa fa_s1_c118_n603 (
        .a(stage1_col118[3]),
        .b(stage1_col118[4]),
        .c_in(stage1_col118[5]),
        .s(fa_s1_c118_n603_s),
        .c_out(fa_s1_c118_n603_c)
    );

    fa fa_s1_c118_n604 (
        .a(stage1_col118[6]),
        .b(stage1_col118[7]),
        .c_in(stage1_col118[8]),
        .s(fa_s1_c118_n604_s),
        .c_out(fa_s1_c118_n604_c)
    );

    fa fa_s1_c118_n605 (
        .a(stage1_col118[9]),
        .b(stage1_col118[10]),
        .c_in(stage1_col118[11]),
        .s(fa_s1_c118_n605_s),
        .c_out(fa_s1_c118_n605_c)
    );

    fa fa_s1_c118_n606 (
        .a(stage1_col118[12]),
        .b(stage1_col118[13]),
        .c_in(stage1_col118[14]),
        .s(fa_s1_c118_n606_s),
        .c_out(fa_s1_c118_n606_c)
    );

    fa fa_s1_c118_n607 (
        .a(stage1_col118[15]),
        .b(stage1_col118[16]),
        .c_in(stage1_col118[17]),
        .s(fa_s1_c118_n607_s),
        .c_out(fa_s1_c118_n607_c)
    );

    fa fa_s1_c118_n608 (
        .a(stage1_col118[18]),
        .b(stage1_col118[19]),
        .c_in(stage1_col118[20]),
        .s(fa_s1_c118_n608_s),
        .c_out(fa_s1_c118_n608_c)
    );

    fa fa_s1_c119_n609 (
        .a(stage1_col119[0]),
        .b(stage1_col119[1]),
        .c_in(stage1_col119[2]),
        .s(fa_s1_c119_n609_s),
        .c_out(fa_s1_c119_n609_c)
    );

    fa fa_s1_c119_n610 (
        .a(stage1_col119[3]),
        .b(stage1_col119[4]),
        .c_in(stage1_col119[5]),
        .s(fa_s1_c119_n610_s),
        .c_out(fa_s1_c119_n610_c)
    );

    fa fa_s1_c119_n611 (
        .a(stage1_col119[6]),
        .b(stage1_col119[7]),
        .c_in(stage1_col119[8]),
        .s(fa_s1_c119_n611_s),
        .c_out(fa_s1_c119_n611_c)
    );

    fa fa_s1_c119_n612 (
        .a(stage1_col119[9]),
        .b(stage1_col119[10]),
        .c_in(stage1_col119[11]),
        .s(fa_s1_c119_n612_s),
        .c_out(fa_s1_c119_n612_c)
    );

    fa fa_s1_c119_n613 (
        .a(stage1_col119[12]),
        .b(stage1_col119[13]),
        .c_in(stage1_col119[14]),
        .s(fa_s1_c119_n613_s),
        .c_out(fa_s1_c119_n613_c)
    );

    fa fa_s1_c119_n614 (
        .a(stage1_col119[15]),
        .b(stage1_col119[16]),
        .c_in(stage1_col119[17]),
        .s(fa_s1_c119_n614_s),
        .c_out(fa_s1_c119_n614_c)
    );

    fa fa_s1_c119_n615 (
        .a(stage1_col119[18]),
        .b(stage1_col119[19]),
        .c_in(stage1_col119[20]),
        .s(fa_s1_c119_n615_s),
        .c_out(fa_s1_c119_n615_c)
    );

    fa fa_s1_c120_n616 (
        .a(stage1_col120[0]),
        .b(stage1_col120[1]),
        .c_in(stage1_col120[2]),
        .s(fa_s1_c120_n616_s),
        .c_out(fa_s1_c120_n616_c)
    );

    fa fa_s1_c120_n617 (
        .a(stage1_col120[3]),
        .b(stage1_col120[4]),
        .c_in(stage1_col120[5]),
        .s(fa_s1_c120_n617_s),
        .c_out(fa_s1_c120_n617_c)
    );

    fa fa_s1_c120_n618 (
        .a(stage1_col120[6]),
        .b(stage1_col120[7]),
        .c_in(stage1_col120[8]),
        .s(fa_s1_c120_n618_s),
        .c_out(fa_s1_c120_n618_c)
    );

    fa fa_s1_c120_n619 (
        .a(stage1_col120[9]),
        .b(stage1_col120[10]),
        .c_in(stage1_col120[11]),
        .s(fa_s1_c120_n619_s),
        .c_out(fa_s1_c120_n619_c)
    );

    fa fa_s1_c120_n620 (
        .a(stage1_col120[12]),
        .b(stage1_col120[13]),
        .c_in(stage1_col120[14]),
        .s(fa_s1_c120_n620_s),
        .c_out(fa_s1_c120_n620_c)
    );

    fa fa_s1_c120_n621 (
        .a(stage1_col120[15]),
        .b(stage1_col120[16]),
        .c_in(stage1_col120[17]),
        .s(fa_s1_c120_n621_s),
        .c_out(fa_s1_c120_n621_c)
    );

    fa fa_s1_c120_n622 (
        .a(stage1_col120[18]),
        .b(stage1_col120[19]),
        .c_in(stage1_col120[20]),
        .s(fa_s1_c120_n622_s),
        .c_out(fa_s1_c120_n622_c)
    );

    fa fa_s1_c121_n623 (
        .a(stage1_col121[0]),
        .b(stage1_col121[1]),
        .c_in(stage1_col121[2]),
        .s(fa_s1_c121_n623_s),
        .c_out(fa_s1_c121_n623_c)
    );

    fa fa_s1_c121_n624 (
        .a(stage1_col121[3]),
        .b(stage1_col121[4]),
        .c_in(stage1_col121[5]),
        .s(fa_s1_c121_n624_s),
        .c_out(fa_s1_c121_n624_c)
    );

    fa fa_s1_c121_n625 (
        .a(stage1_col121[6]),
        .b(stage1_col121[7]),
        .c_in(stage1_col121[8]),
        .s(fa_s1_c121_n625_s),
        .c_out(fa_s1_c121_n625_c)
    );

    fa fa_s1_c121_n626 (
        .a(stage1_col121[9]),
        .b(stage1_col121[10]),
        .c_in(stage1_col121[11]),
        .s(fa_s1_c121_n626_s),
        .c_out(fa_s1_c121_n626_c)
    );

    fa fa_s1_c121_n627 (
        .a(stage1_col121[12]),
        .b(stage1_col121[13]),
        .c_in(stage1_col121[14]),
        .s(fa_s1_c121_n627_s),
        .c_out(fa_s1_c121_n627_c)
    );

    fa fa_s1_c121_n628 (
        .a(stage1_col121[15]),
        .b(stage1_col121[16]),
        .c_in(stage1_col121[17]),
        .s(fa_s1_c121_n628_s),
        .c_out(fa_s1_c121_n628_c)
    );

    fa fa_s1_c121_n629 (
        .a(stage1_col121[18]),
        .b(stage1_col121[19]),
        .c_in(stage1_col121[20]),
        .s(fa_s1_c121_n629_s),
        .c_out(fa_s1_c121_n629_c)
    );

    fa fa_s1_c122_n630 (
        .a(stage1_col122[0]),
        .b(stage1_col122[1]),
        .c_in(stage1_col122[2]),
        .s(fa_s1_c122_n630_s),
        .c_out(fa_s1_c122_n630_c)
    );

    fa fa_s1_c122_n631 (
        .a(stage1_col122[3]),
        .b(stage1_col122[4]),
        .c_in(stage1_col122[5]),
        .s(fa_s1_c122_n631_s),
        .c_out(fa_s1_c122_n631_c)
    );

    fa fa_s1_c122_n632 (
        .a(stage1_col122[6]),
        .b(stage1_col122[7]),
        .c_in(stage1_col122[8]),
        .s(fa_s1_c122_n632_s),
        .c_out(fa_s1_c122_n632_c)
    );

    fa fa_s1_c122_n633 (
        .a(stage1_col122[9]),
        .b(stage1_col122[10]),
        .c_in(stage1_col122[11]),
        .s(fa_s1_c122_n633_s),
        .c_out(fa_s1_c122_n633_c)
    );

    fa fa_s1_c122_n634 (
        .a(stage1_col122[12]),
        .b(stage1_col122[13]),
        .c_in(stage1_col122[14]),
        .s(fa_s1_c122_n634_s),
        .c_out(fa_s1_c122_n634_c)
    );

    fa fa_s1_c122_n635 (
        .a(stage1_col122[15]),
        .b(stage1_col122[16]),
        .c_in(stage1_col122[17]),
        .s(fa_s1_c122_n635_s),
        .c_out(fa_s1_c122_n635_c)
    );

    fa fa_s1_c122_n636 (
        .a(stage1_col122[18]),
        .b(stage1_col122[19]),
        .c_in(stage1_col122[20]),
        .s(fa_s1_c122_n636_s),
        .c_out(fa_s1_c122_n636_c)
    );

    fa fa_s1_c123_n637 (
        .a(stage1_col123[0]),
        .b(stage1_col123[1]),
        .c_in(stage1_col123[2]),
        .s(fa_s1_c123_n637_s),
        .c_out(fa_s1_c123_n637_c)
    );

    fa fa_s1_c123_n638 (
        .a(stage1_col123[3]),
        .b(stage1_col123[4]),
        .c_in(stage1_col123[5]),
        .s(fa_s1_c123_n638_s),
        .c_out(fa_s1_c123_n638_c)
    );

    fa fa_s1_c123_n639 (
        .a(stage1_col123[6]),
        .b(stage1_col123[7]),
        .c_in(stage1_col123[8]),
        .s(fa_s1_c123_n639_s),
        .c_out(fa_s1_c123_n639_c)
    );

    fa fa_s1_c123_n640 (
        .a(stage1_col123[9]),
        .b(stage1_col123[10]),
        .c_in(stage1_col123[11]),
        .s(fa_s1_c123_n640_s),
        .c_out(fa_s1_c123_n640_c)
    );

    fa fa_s1_c123_n641 (
        .a(stage1_col123[12]),
        .b(stage1_col123[13]),
        .c_in(stage1_col123[14]),
        .s(fa_s1_c123_n641_s),
        .c_out(fa_s1_c123_n641_c)
    );

    fa fa_s1_c123_n642 (
        .a(stage1_col123[15]),
        .b(stage1_col123[16]),
        .c_in(stage1_col123[17]),
        .s(fa_s1_c123_n642_s),
        .c_out(fa_s1_c123_n642_c)
    );

    fa fa_s1_c123_n643 (
        .a(stage1_col123[18]),
        .b(stage1_col123[19]),
        .c_in(stage1_col123[20]),
        .s(fa_s1_c123_n643_s),
        .c_out(fa_s1_c123_n643_c)
    );

    fa fa_s1_c124_n644 (
        .a(stage1_col124[0]),
        .b(stage1_col124[1]),
        .c_in(stage1_col124[2]),
        .s(fa_s1_c124_n644_s),
        .c_out(fa_s1_c124_n644_c)
    );

    fa fa_s1_c124_n645 (
        .a(stage1_col124[3]),
        .b(stage1_col124[4]),
        .c_in(stage1_col124[5]),
        .s(fa_s1_c124_n645_s),
        .c_out(fa_s1_c124_n645_c)
    );

    fa fa_s1_c124_n646 (
        .a(stage1_col124[6]),
        .b(stage1_col124[7]),
        .c_in(stage1_col124[8]),
        .s(fa_s1_c124_n646_s),
        .c_out(fa_s1_c124_n646_c)
    );

    fa fa_s1_c124_n647 (
        .a(stage1_col124[9]),
        .b(stage1_col124[10]),
        .c_in(stage1_col124[11]),
        .s(fa_s1_c124_n647_s),
        .c_out(fa_s1_c124_n647_c)
    );

    fa fa_s1_c124_n648 (
        .a(stage1_col124[12]),
        .b(stage1_col124[13]),
        .c_in(stage1_col124[14]),
        .s(fa_s1_c124_n648_s),
        .c_out(fa_s1_c124_n648_c)
    );

    fa fa_s1_c124_n649 (
        .a(stage1_col124[15]),
        .b(stage1_col124[16]),
        .c_in(stage1_col124[17]),
        .s(fa_s1_c124_n649_s),
        .c_out(fa_s1_c124_n649_c)
    );

    fa fa_s1_c124_n650 (
        .a(stage1_col124[18]),
        .b(stage1_col124[19]),
        .c_in(stage1_col124[20]),
        .s(fa_s1_c124_n650_s),
        .c_out(fa_s1_c124_n650_c)
    );

    fa fa_s1_c125_n651 (
        .a(stage1_col125[0]),
        .b(stage1_col125[1]),
        .c_in(stage1_col125[2]),
        .s(fa_s1_c125_n651_s),
        .c_out(fa_s1_c125_n651_c)
    );

    fa fa_s1_c125_n652 (
        .a(stage1_col125[3]),
        .b(stage1_col125[4]),
        .c_in(stage1_col125[5]),
        .s(fa_s1_c125_n652_s),
        .c_out(fa_s1_c125_n652_c)
    );

    fa fa_s1_c125_n653 (
        .a(stage1_col125[6]),
        .b(stage1_col125[7]),
        .c_in(stage1_col125[8]),
        .s(fa_s1_c125_n653_s),
        .c_out(fa_s1_c125_n653_c)
    );

    fa fa_s1_c125_n654 (
        .a(stage1_col125[9]),
        .b(stage1_col125[10]),
        .c_in(stage1_col125[11]),
        .s(fa_s1_c125_n654_s),
        .c_out(fa_s1_c125_n654_c)
    );

    fa fa_s1_c125_n655 (
        .a(stage1_col125[12]),
        .b(stage1_col125[13]),
        .c_in(stage1_col125[14]),
        .s(fa_s1_c125_n655_s),
        .c_out(fa_s1_c125_n655_c)
    );

    fa fa_s1_c125_n656 (
        .a(stage1_col125[15]),
        .b(stage1_col125[16]),
        .c_in(stage1_col125[17]),
        .s(fa_s1_c125_n656_s),
        .c_out(fa_s1_c125_n656_c)
    );

    fa fa_s1_c125_n657 (
        .a(stage1_col125[18]),
        .b(stage1_col125[19]),
        .c_in(stage1_col125[20]),
        .s(fa_s1_c125_n657_s),
        .c_out(fa_s1_c125_n657_c)
    );

    fa fa_s1_c126_n658 (
        .a(stage1_col126[0]),
        .b(stage1_col126[1]),
        .c_in(stage1_col126[2]),
        .s(fa_s1_c126_n658_s),
        .c_out(fa_s1_c126_n658_c)
    );

    fa fa_s1_c126_n659 (
        .a(stage1_col126[3]),
        .b(stage1_col126[4]),
        .c_in(stage1_col126[5]),
        .s(fa_s1_c126_n659_s),
        .c_out(fa_s1_c126_n659_c)
    );

    fa fa_s1_c126_n660 (
        .a(stage1_col126[6]),
        .b(stage1_col126[7]),
        .c_in(stage1_col126[8]),
        .s(fa_s1_c126_n660_s),
        .c_out(fa_s1_c126_n660_c)
    );

    fa fa_s1_c126_n661 (
        .a(stage1_col126[9]),
        .b(stage1_col126[10]),
        .c_in(stage1_col126[11]),
        .s(fa_s1_c126_n661_s),
        .c_out(fa_s1_c126_n661_c)
    );

    fa fa_s1_c126_n662 (
        .a(stage1_col126[12]),
        .b(stage1_col126[13]),
        .c_in(stage1_col126[14]),
        .s(fa_s1_c126_n662_s),
        .c_out(fa_s1_c126_n662_c)
    );

    fa fa_s1_c126_n663 (
        .a(stage1_col126[15]),
        .b(stage1_col126[16]),
        .c_in(stage1_col126[17]),
        .s(fa_s1_c126_n663_s),
        .c_out(fa_s1_c126_n663_c)
    );

    fa fa_s1_c126_n664 (
        .a(stage1_col126[18]),
        .b(stage1_col126[19]),
        .c_in(stage1_col126[20]),
        .s(fa_s1_c126_n664_s),
        .c_out(fa_s1_c126_n664_c)
    );

    ha ha_s1_c1_n0 (
        .a(stage1_col1[0]),
        .b(stage1_col1[1]),
        .s(ha_s1_c1_n0_s),
        .c_out(ha_s1_c1_n0_c)
    );

    // Map to Stage 2 columns
    generate
        if (PIPE) begin : gen_stage2_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage2_col0[0] <= 1'b0;
                    stage2_col1[0] <= 1'b0;
                    stage2_col2[0] <= 1'b0;
                    stage2_col2[1] <= 1'b0;
                    stage2_col3[0] <= 1'b0;
                    stage2_col4[0] <= 1'b0;
                    stage2_col4[1] <= 1'b0;
                    stage2_col4[2] <= 1'b0;
                    stage2_col5[0] <= 1'b0;
                    stage2_col5[1] <= 1'b0;
                    stage2_col6[0] <= 1'b0;
                    stage2_col6[1] <= 1'b0;
                    stage2_col7[0] <= 1'b0;
                    stage2_col7[1] <= 1'b0;
                    stage2_col8[0] <= 1'b0;
                    stage2_col8[1] <= 1'b0;
                    stage2_col9[0] <= 1'b0;
                    stage2_col9[1] <= 1'b0;
                    stage2_col9[2] <= 1'b0;
                    stage2_col9[3] <= 1'b0;
                    stage2_col10[0] <= 1'b0;
                    stage2_col10[1] <= 1'b0;
                    stage2_col10[2] <= 1'b0;
                    stage2_col11[0] <= 1'b0;
                    stage2_col11[1] <= 1'b0;
                    stage2_col11[2] <= 1'b0;
                    stage2_col12[0] <= 1'b0;
                    stage2_col12[1] <= 1'b0;
                    stage2_col12[2] <= 1'b0;
                    stage2_col13[0] <= 1'b0;
                    stage2_col13[1] <= 1'b0;
                    stage2_col13[2] <= 1'b0;
                    stage2_col13[3] <= 1'b0;
                    stage2_col13[4] <= 1'b0;
                    stage2_col14[0] <= 1'b0;
                    stage2_col14[1] <= 1'b0;
                    stage2_col14[2] <= 1'b0;
                    stage2_col14[3] <= 1'b0;
                    stage2_col15[0] <= 1'b0;
                    stage2_col15[1] <= 1'b0;
                    stage2_col15[2] <= 1'b0;
                    stage2_col15[3] <= 1'b0;
                    stage2_col16[0] <= 1'b0;
                    stage2_col16[1] <= 1'b0;
                    stage2_col16[2] <= 1'b0;
                    stage2_col16[3] <= 1'b0;
                    stage2_col17[0] <= 1'b0;
                    stage2_col17[1] <= 1'b0;
                    stage2_col17[2] <= 1'b0;
                    stage2_col17[3] <= 1'b0;
                    stage2_col18[0] <= 1'b0;
                    stage2_col18[1] <= 1'b0;
                    stage2_col18[2] <= 1'b0;
                    stage2_col18[3] <= 1'b0;
                    stage2_col18[4] <= 1'b0;
                    stage2_col18[5] <= 1'b0;
                    stage2_col19[0] <= 1'b0;
                    stage2_col19[1] <= 1'b0;
                    stage2_col19[2] <= 1'b0;
                    stage2_col19[3] <= 1'b0;
                    stage2_col19[4] <= 1'b0;
                    stage2_col20[0] <= 1'b0;
                    stage2_col20[1] <= 1'b0;
                    stage2_col20[2] <= 1'b0;
                    stage2_col20[3] <= 1'b0;
                    stage2_col20[4] <= 1'b0;
                    stage2_col21[0] <= 1'b0;
                    stage2_col21[1] <= 1'b0;
                    stage2_col21[2] <= 1'b0;
                    stage2_col21[3] <= 1'b0;
                    stage2_col21[4] <= 1'b0;
                    stage2_col22[0] <= 1'b0;
                    stage2_col22[1] <= 1'b0;
                    stage2_col22[2] <= 1'b0;
                    stage2_col22[3] <= 1'b0;
                    stage2_col22[4] <= 1'b0;
                    stage2_col22[5] <= 1'b0;
                    stage2_col22[6] <= 1'b0;
                    stage2_col23[0] <= 1'b0;
                    stage2_col23[1] <= 1'b0;
                    stage2_col23[2] <= 1'b0;
                    stage2_col23[3] <= 1'b0;
                    stage2_col23[4] <= 1'b0;
                    stage2_col23[5] <= 1'b0;
                    stage2_col24[0] <= 1'b0;
                    stage2_col24[1] <= 1'b0;
                    stage2_col24[2] <= 1'b0;
                    stage2_col24[3] <= 1'b0;
                    stage2_col24[4] <= 1'b0;
                    stage2_col24[5] <= 1'b0;
                    stage2_col25[0] <= 1'b0;
                    stage2_col25[1] <= 1'b0;
                    stage2_col25[2] <= 1'b0;
                    stage2_col25[3] <= 1'b0;
                    stage2_col25[4] <= 1'b0;
                    stage2_col25[5] <= 1'b0;
                    stage2_col26[0] <= 1'b0;
                    stage2_col26[1] <= 1'b0;
                    stage2_col26[2] <= 1'b0;
                    stage2_col26[3] <= 1'b0;
                    stage2_col26[4] <= 1'b0;
                    stage2_col26[5] <= 1'b0;
                    stage2_col27[0] <= 1'b0;
                    stage2_col27[1] <= 1'b0;
                    stage2_col27[2] <= 1'b0;
                    stage2_col27[3] <= 1'b0;
                    stage2_col27[4] <= 1'b0;
                    stage2_col27[5] <= 1'b0;
                    stage2_col27[6] <= 1'b0;
                    stage2_col27[7] <= 1'b0;
                    stage2_col28[0] <= 1'b0;
                    stage2_col28[1] <= 1'b0;
                    stage2_col28[2] <= 1'b0;
                    stage2_col28[3] <= 1'b0;
                    stage2_col28[4] <= 1'b0;
                    stage2_col28[5] <= 1'b0;
                    stage2_col28[6] <= 1'b0;
                    stage2_col29[0] <= 1'b0;
                    stage2_col29[1] <= 1'b0;
                    stage2_col29[2] <= 1'b0;
                    stage2_col29[3] <= 1'b0;
                    stage2_col29[4] <= 1'b0;
                    stage2_col29[5] <= 1'b0;
                    stage2_col29[6] <= 1'b0;
                    stage2_col30[0] <= 1'b0;
                    stage2_col30[1] <= 1'b0;
                    stage2_col30[2] <= 1'b0;
                    stage2_col30[3] <= 1'b0;
                    stage2_col30[4] <= 1'b0;
                    stage2_col30[5] <= 1'b0;
                    stage2_col30[6] <= 1'b0;
                    stage2_col31[0] <= 1'b0;
                    stage2_col31[1] <= 1'b0;
                    stage2_col31[2] <= 1'b0;
                    stage2_col31[3] <= 1'b0;
                    stage2_col31[4] <= 1'b0;
                    stage2_col31[5] <= 1'b0;
                    stage2_col31[6] <= 1'b0;
                    stage2_col31[7] <= 1'b0;
                    stage2_col31[8] <= 1'b0;
                    stage2_col32[0] <= 1'b0;
                    stage2_col32[1] <= 1'b0;
                    stage2_col32[2] <= 1'b0;
                    stage2_col32[3] <= 1'b0;
                    stage2_col32[4] <= 1'b0;
                    stage2_col32[5] <= 1'b0;
                    stage2_col32[6] <= 1'b0;
                    stage2_col32[7] <= 1'b0;
                    stage2_col33[0] <= 1'b0;
                    stage2_col33[1] <= 1'b0;
                    stage2_col33[2] <= 1'b0;
                    stage2_col33[3] <= 1'b0;
                    stage2_col33[4] <= 1'b0;
                    stage2_col33[5] <= 1'b0;
                    stage2_col33[6] <= 1'b0;
                    stage2_col33[7] <= 1'b0;
                    stage2_col34[0] <= 1'b0;
                    stage2_col34[1] <= 1'b0;
                    stage2_col34[2] <= 1'b0;
                    stage2_col34[3] <= 1'b0;
                    stage2_col34[4] <= 1'b0;
                    stage2_col34[5] <= 1'b0;
                    stage2_col34[6] <= 1'b0;
                    stage2_col34[7] <= 1'b0;
                    stage2_col35[0] <= 1'b0;
                    stage2_col35[1] <= 1'b0;
                    stage2_col35[2] <= 1'b0;
                    stage2_col35[3] <= 1'b0;
                    stage2_col35[4] <= 1'b0;
                    stage2_col35[5] <= 1'b0;
                    stage2_col35[6] <= 1'b0;
                    stage2_col35[7] <= 1'b0;
                    stage2_col36[0] <= 1'b0;
                    stage2_col36[1] <= 1'b0;
                    stage2_col36[2] <= 1'b0;
                    stage2_col36[3] <= 1'b0;
                    stage2_col36[4] <= 1'b0;
                    stage2_col36[5] <= 1'b0;
                    stage2_col36[6] <= 1'b0;
                    stage2_col36[7] <= 1'b0;
                    stage2_col36[8] <= 1'b0;
                    stage2_col36[9] <= 1'b0;
                    stage2_col37[0] <= 1'b0;
                    stage2_col37[1] <= 1'b0;
                    stage2_col37[2] <= 1'b0;
                    stage2_col37[3] <= 1'b0;
                    stage2_col37[4] <= 1'b0;
                    stage2_col37[5] <= 1'b0;
                    stage2_col37[6] <= 1'b0;
                    stage2_col37[7] <= 1'b0;
                    stage2_col37[8] <= 1'b0;
                    stage2_col38[0] <= 1'b0;
                    stage2_col38[1] <= 1'b0;
                    stage2_col38[2] <= 1'b0;
                    stage2_col38[3] <= 1'b0;
                    stage2_col38[4] <= 1'b0;
                    stage2_col38[5] <= 1'b0;
                    stage2_col38[6] <= 1'b0;
                    stage2_col38[7] <= 1'b0;
                    stage2_col38[8] <= 1'b0;
                    stage2_col39[0] <= 1'b0;
                    stage2_col39[1] <= 1'b0;
                    stage2_col39[2] <= 1'b0;
                    stage2_col39[3] <= 1'b0;
                    stage2_col39[4] <= 1'b0;
                    stage2_col39[5] <= 1'b0;
                    stage2_col39[6] <= 1'b0;
                    stage2_col39[7] <= 1'b0;
                    stage2_col39[8] <= 1'b0;
                    stage2_col40[0] <= 1'b0;
                    stage2_col40[1] <= 1'b0;
                    stage2_col40[2] <= 1'b0;
                    stage2_col40[3] <= 1'b0;
                    stage2_col40[4] <= 1'b0;
                    stage2_col40[5] <= 1'b0;
                    stage2_col40[6] <= 1'b0;
                    stage2_col40[7] <= 1'b0;
                    stage2_col40[8] <= 1'b0;
                    stage2_col40[9] <= 1'b0;
                    stage2_col40[10] <= 1'b0;
                    stage2_col41[0] <= 1'b0;
                    stage2_col41[1] <= 1'b0;
                    stage2_col41[2] <= 1'b0;
                    stage2_col41[3] <= 1'b0;
                    stage2_col41[4] <= 1'b0;
                    stage2_col41[5] <= 1'b0;
                    stage2_col41[6] <= 1'b0;
                    stage2_col41[7] <= 1'b0;
                    stage2_col41[8] <= 1'b0;
                    stage2_col41[9] <= 1'b0;
                    stage2_col42[0] <= 1'b0;
                    stage2_col42[1] <= 1'b0;
                    stage2_col42[2] <= 1'b0;
                    stage2_col42[3] <= 1'b0;
                    stage2_col42[4] <= 1'b0;
                    stage2_col42[5] <= 1'b0;
                    stage2_col42[6] <= 1'b0;
                    stage2_col42[7] <= 1'b0;
                    stage2_col42[8] <= 1'b0;
                    stage2_col42[9] <= 1'b0;
                    stage2_col43[0] <= 1'b0;
                    stage2_col43[1] <= 1'b0;
                    stage2_col43[2] <= 1'b0;
                    stage2_col43[3] <= 1'b0;
                    stage2_col43[4] <= 1'b0;
                    stage2_col43[5] <= 1'b0;
                    stage2_col43[6] <= 1'b0;
                    stage2_col43[7] <= 1'b0;
                    stage2_col43[8] <= 1'b0;
                    stage2_col43[9] <= 1'b0;
                    stage2_col44[0] <= 1'b0;
                    stage2_col44[1] <= 1'b0;
                    stage2_col44[2] <= 1'b0;
                    stage2_col44[3] <= 1'b0;
                    stage2_col44[4] <= 1'b0;
                    stage2_col44[5] <= 1'b0;
                    stage2_col44[6] <= 1'b0;
                    stage2_col44[7] <= 1'b0;
                    stage2_col44[8] <= 1'b0;
                    stage2_col44[9] <= 1'b0;
                    stage2_col45[0] <= 1'b0;
                    stage2_col45[1] <= 1'b0;
                    stage2_col45[2] <= 1'b0;
                    stage2_col45[3] <= 1'b0;
                    stage2_col45[4] <= 1'b0;
                    stage2_col45[5] <= 1'b0;
                    stage2_col45[6] <= 1'b0;
                    stage2_col45[7] <= 1'b0;
                    stage2_col45[8] <= 1'b0;
                    stage2_col45[9] <= 1'b0;
                    stage2_col45[10] <= 1'b0;
                    stage2_col45[11] <= 1'b0;
                    stage2_col46[0] <= 1'b0;
                    stage2_col46[1] <= 1'b0;
                    stage2_col46[2] <= 1'b0;
                    stage2_col46[3] <= 1'b0;
                    stage2_col46[4] <= 1'b0;
                    stage2_col46[5] <= 1'b0;
                    stage2_col46[6] <= 1'b0;
                    stage2_col46[7] <= 1'b0;
                    stage2_col46[8] <= 1'b0;
                    stage2_col46[9] <= 1'b0;
                    stage2_col46[10] <= 1'b0;
                    stage2_col47[0] <= 1'b0;
                    stage2_col47[1] <= 1'b0;
                    stage2_col47[2] <= 1'b0;
                    stage2_col47[3] <= 1'b0;
                    stage2_col47[4] <= 1'b0;
                    stage2_col47[5] <= 1'b0;
                    stage2_col47[6] <= 1'b0;
                    stage2_col47[7] <= 1'b0;
                    stage2_col47[8] <= 1'b0;
                    stage2_col47[9] <= 1'b0;
                    stage2_col47[10] <= 1'b0;
                    stage2_col48[0] <= 1'b0;
                    stage2_col48[1] <= 1'b0;
                    stage2_col48[2] <= 1'b0;
                    stage2_col48[3] <= 1'b0;
                    stage2_col48[4] <= 1'b0;
                    stage2_col48[5] <= 1'b0;
                    stage2_col48[6] <= 1'b0;
                    stage2_col48[7] <= 1'b0;
                    stage2_col48[8] <= 1'b0;
                    stage2_col48[9] <= 1'b0;
                    stage2_col48[10] <= 1'b0;
                    stage2_col49[0] <= 1'b0;
                    stage2_col49[1] <= 1'b0;
                    stage2_col49[2] <= 1'b0;
                    stage2_col49[3] <= 1'b0;
                    stage2_col49[4] <= 1'b0;
                    stage2_col49[5] <= 1'b0;
                    stage2_col49[6] <= 1'b0;
                    stage2_col49[7] <= 1'b0;
                    stage2_col49[8] <= 1'b0;
                    stage2_col49[9] <= 1'b0;
                    stage2_col49[10] <= 1'b0;
                    stage2_col49[11] <= 1'b0;
                    stage2_col49[12] <= 1'b0;
                    stage2_col50[0] <= 1'b0;
                    stage2_col50[1] <= 1'b0;
                    stage2_col50[2] <= 1'b0;
                    stage2_col50[3] <= 1'b0;
                    stage2_col50[4] <= 1'b0;
                    stage2_col50[5] <= 1'b0;
                    stage2_col50[6] <= 1'b0;
                    stage2_col50[7] <= 1'b0;
                    stage2_col50[8] <= 1'b0;
                    stage2_col50[9] <= 1'b0;
                    stage2_col50[10] <= 1'b0;
                    stage2_col50[11] <= 1'b0;
                    stage2_col51[0] <= 1'b0;
                    stage2_col51[1] <= 1'b0;
                    stage2_col51[2] <= 1'b0;
                    stage2_col51[3] <= 1'b0;
                    stage2_col51[4] <= 1'b0;
                    stage2_col51[5] <= 1'b0;
                    stage2_col51[6] <= 1'b0;
                    stage2_col51[7] <= 1'b0;
                    stage2_col51[8] <= 1'b0;
                    stage2_col51[9] <= 1'b0;
                    stage2_col51[10] <= 1'b0;
                    stage2_col51[11] <= 1'b0;
                    stage2_col52[0] <= 1'b0;
                    stage2_col52[1] <= 1'b0;
                    stage2_col52[2] <= 1'b0;
                    stage2_col52[3] <= 1'b0;
                    stage2_col52[4] <= 1'b0;
                    stage2_col52[5] <= 1'b0;
                    stage2_col52[6] <= 1'b0;
                    stage2_col52[7] <= 1'b0;
                    stage2_col52[8] <= 1'b0;
                    stage2_col52[9] <= 1'b0;
                    stage2_col52[10] <= 1'b0;
                    stage2_col52[11] <= 1'b0;
                    stage2_col53[0] <= 1'b0;
                    stage2_col53[1] <= 1'b0;
                    stage2_col53[2] <= 1'b0;
                    stage2_col53[3] <= 1'b0;
                    stage2_col53[4] <= 1'b0;
                    stage2_col53[5] <= 1'b0;
                    stage2_col53[6] <= 1'b0;
                    stage2_col53[7] <= 1'b0;
                    stage2_col53[8] <= 1'b0;
                    stage2_col53[9] <= 1'b0;
                    stage2_col53[10] <= 1'b0;
                    stage2_col53[11] <= 1'b0;
                    stage2_col54[0] <= 1'b0;
                    stage2_col54[1] <= 1'b0;
                    stage2_col54[2] <= 1'b0;
                    stage2_col54[3] <= 1'b0;
                    stage2_col54[4] <= 1'b0;
                    stage2_col54[5] <= 1'b0;
                    stage2_col54[6] <= 1'b0;
                    stage2_col54[7] <= 1'b0;
                    stage2_col54[8] <= 1'b0;
                    stage2_col54[9] <= 1'b0;
                    stage2_col54[10] <= 1'b0;
                    stage2_col54[11] <= 1'b0;
                    stage2_col54[12] <= 1'b0;
                    stage2_col54[13] <= 1'b0;
                    stage2_col55[0] <= 1'b0;
                    stage2_col55[1] <= 1'b0;
                    stage2_col55[2] <= 1'b0;
                    stage2_col55[3] <= 1'b0;
                    stage2_col55[4] <= 1'b0;
                    stage2_col55[5] <= 1'b0;
                    stage2_col55[6] <= 1'b0;
                    stage2_col55[7] <= 1'b0;
                    stage2_col55[8] <= 1'b0;
                    stage2_col55[9] <= 1'b0;
                    stage2_col55[10] <= 1'b0;
                    stage2_col55[11] <= 1'b0;
                    stage2_col55[12] <= 1'b0;
                    stage2_col56[0] <= 1'b0;
                    stage2_col56[1] <= 1'b0;
                    stage2_col56[2] <= 1'b0;
                    stage2_col56[3] <= 1'b0;
                    stage2_col56[4] <= 1'b0;
                    stage2_col56[5] <= 1'b0;
                    stage2_col56[6] <= 1'b0;
                    stage2_col56[7] <= 1'b0;
                    stage2_col56[8] <= 1'b0;
                    stage2_col56[9] <= 1'b0;
                    stage2_col56[10] <= 1'b0;
                    stage2_col56[11] <= 1'b0;
                    stage2_col56[12] <= 1'b0;
                    stage2_col57[0] <= 1'b0;
                    stage2_col57[1] <= 1'b0;
                    stage2_col57[2] <= 1'b0;
                    stage2_col57[3] <= 1'b0;
                    stage2_col57[4] <= 1'b0;
                    stage2_col57[5] <= 1'b0;
                    stage2_col57[6] <= 1'b0;
                    stage2_col57[7] <= 1'b0;
                    stage2_col57[8] <= 1'b0;
                    stage2_col57[9] <= 1'b0;
                    stage2_col57[10] <= 1'b0;
                    stage2_col57[11] <= 1'b0;
                    stage2_col57[12] <= 1'b0;
                    stage2_col58[0] <= 1'b0;
                    stage2_col58[1] <= 1'b0;
                    stage2_col58[2] <= 1'b0;
                    stage2_col58[3] <= 1'b0;
                    stage2_col58[4] <= 1'b0;
                    stage2_col58[5] <= 1'b0;
                    stage2_col58[6] <= 1'b0;
                    stage2_col58[7] <= 1'b0;
                    stage2_col58[8] <= 1'b0;
                    stage2_col58[9] <= 1'b0;
                    stage2_col58[10] <= 1'b0;
                    stage2_col58[11] <= 1'b0;
                    stage2_col58[12] <= 1'b0;
                    stage2_col58[13] <= 1'b0;
                    stage2_col58[14] <= 1'b0;
                    stage2_col59[0] <= 1'b0;
                    stage2_col59[1] <= 1'b0;
                    stage2_col59[2] <= 1'b0;
                    stage2_col59[3] <= 1'b0;
                    stage2_col59[4] <= 1'b0;
                    stage2_col59[5] <= 1'b0;
                    stage2_col59[6] <= 1'b0;
                    stage2_col59[7] <= 1'b0;
                    stage2_col59[8] <= 1'b0;
                    stage2_col59[9] <= 1'b0;
                    stage2_col59[10] <= 1'b0;
                    stage2_col59[11] <= 1'b0;
                    stage2_col59[12] <= 1'b0;
                    stage2_col59[13] <= 1'b0;
                    stage2_col60[0] <= 1'b0;
                    stage2_col60[1] <= 1'b0;
                    stage2_col60[2] <= 1'b0;
                    stage2_col60[3] <= 1'b0;
                    stage2_col60[4] <= 1'b0;
                    stage2_col60[5] <= 1'b0;
                    stage2_col60[6] <= 1'b0;
                    stage2_col60[7] <= 1'b0;
                    stage2_col60[8] <= 1'b0;
                    stage2_col60[9] <= 1'b0;
                    stage2_col60[10] <= 1'b0;
                    stage2_col60[11] <= 1'b0;
                    stage2_col60[12] <= 1'b0;
                    stage2_col60[13] <= 1'b0;
                    stage2_col61[0] <= 1'b0;
                    stage2_col61[1] <= 1'b0;
                    stage2_col61[2] <= 1'b0;
                    stage2_col61[3] <= 1'b0;
                    stage2_col61[4] <= 1'b0;
                    stage2_col61[5] <= 1'b0;
                    stage2_col61[6] <= 1'b0;
                    stage2_col61[7] <= 1'b0;
                    stage2_col61[8] <= 1'b0;
                    stage2_col61[9] <= 1'b0;
                    stage2_col61[10] <= 1'b0;
                    stage2_col61[11] <= 1'b0;
                    stage2_col61[12] <= 1'b0;
                    stage2_col61[13] <= 1'b0;
                    stage2_col62[0] <= 1'b0;
                    stage2_col62[1] <= 1'b0;
                    stage2_col62[2] <= 1'b0;
                    stage2_col62[3] <= 1'b0;
                    stage2_col62[4] <= 1'b0;
                    stage2_col62[5] <= 1'b0;
                    stage2_col62[6] <= 1'b0;
                    stage2_col62[7] <= 1'b0;
                    stage2_col62[8] <= 1'b0;
                    stage2_col62[9] <= 1'b0;
                    stage2_col62[10] <= 1'b0;
                    stage2_col62[11] <= 1'b0;
                    stage2_col62[12] <= 1'b0;
                    stage2_col62[13] <= 1'b0;
                    stage2_col63[0] <= 1'b0;
                    stage2_col63[1] <= 1'b0;
                    stage2_col63[2] <= 1'b0;
                    stage2_col63[3] <= 1'b0;
                    stage2_col63[4] <= 1'b0;
                    stage2_col63[5] <= 1'b0;
                    stage2_col63[6] <= 1'b0;
                    stage2_col63[7] <= 1'b0;
                    stage2_col63[8] <= 1'b0;
                    stage2_col63[9] <= 1'b0;
                    stage2_col63[10] <= 1'b0;
                    stage2_col63[11] <= 1'b0;
                    stage2_col63[12] <= 1'b0;
                    stage2_col63[13] <= 1'b0;
                    stage2_col63[14] <= 1'b0;
                    stage2_col63[15] <= 1'b0;
                    stage2_col64[0] <= 1'b0;
                    stage2_col64[1] <= 1'b0;
                    stage2_col64[2] <= 1'b0;
                    stage2_col64[3] <= 1'b0;
                    stage2_col64[4] <= 1'b0;
                    stage2_col64[5] <= 1'b0;
                    stage2_col64[6] <= 1'b0;
                    stage2_col64[7] <= 1'b0;
                    stage2_col64[8] <= 1'b0;
                    stage2_col64[9] <= 1'b0;
                    stage2_col64[10] <= 1'b0;
                    stage2_col64[11] <= 1'b0;
                    stage2_col64[12] <= 1'b0;
                    stage2_col64[13] <= 1'b0;
                    stage2_col65[0] <= 1'b0;
                    stage2_col65[1] <= 1'b0;
                    stage2_col65[2] <= 1'b0;
                    stage2_col65[3] <= 1'b0;
                    stage2_col65[4] <= 1'b0;
                    stage2_col65[5] <= 1'b0;
                    stage2_col65[6] <= 1'b0;
                    stage2_col65[7] <= 1'b0;
                    stage2_col65[8] <= 1'b0;
                    stage2_col65[9] <= 1'b0;
                    stage2_col65[10] <= 1'b0;
                    stage2_col65[11] <= 1'b0;
                    stage2_col65[12] <= 1'b0;
                    stage2_col65[13] <= 1'b0;
                    stage2_col65[14] <= 1'b0;
                    stage2_col65[15] <= 1'b0;
                    stage2_col66[0] <= 1'b0;
                    stage2_col66[1] <= 1'b0;
                    stage2_col66[2] <= 1'b0;
                    stage2_col66[3] <= 1'b0;
                    stage2_col66[4] <= 1'b0;
                    stage2_col66[5] <= 1'b0;
                    stage2_col66[6] <= 1'b0;
                    stage2_col66[7] <= 1'b0;
                    stage2_col66[8] <= 1'b0;
                    stage2_col66[9] <= 1'b0;
                    stage2_col66[10] <= 1'b0;
                    stage2_col66[11] <= 1'b0;
                    stage2_col66[12] <= 1'b0;
                    stage2_col66[13] <= 1'b0;
                    stage2_col67[0] <= 1'b0;
                    stage2_col67[1] <= 1'b0;
                    stage2_col67[2] <= 1'b0;
                    stage2_col67[3] <= 1'b0;
                    stage2_col67[4] <= 1'b0;
                    stage2_col67[5] <= 1'b0;
                    stage2_col67[6] <= 1'b0;
                    stage2_col67[7] <= 1'b0;
                    stage2_col67[8] <= 1'b0;
                    stage2_col67[9] <= 1'b0;
                    stage2_col67[10] <= 1'b0;
                    stage2_col67[11] <= 1'b0;
                    stage2_col67[12] <= 1'b0;
                    stage2_col67[13] <= 1'b0;
                    stage2_col67[14] <= 1'b0;
                    stage2_col67[15] <= 1'b0;
                    stage2_col68[0] <= 1'b0;
                    stage2_col68[1] <= 1'b0;
                    stage2_col68[2] <= 1'b0;
                    stage2_col68[3] <= 1'b0;
                    stage2_col68[4] <= 1'b0;
                    stage2_col68[5] <= 1'b0;
                    stage2_col68[6] <= 1'b0;
                    stage2_col68[7] <= 1'b0;
                    stage2_col68[8] <= 1'b0;
                    stage2_col68[9] <= 1'b0;
                    stage2_col68[10] <= 1'b0;
                    stage2_col68[11] <= 1'b0;
                    stage2_col68[12] <= 1'b0;
                    stage2_col68[13] <= 1'b0;
                    stage2_col69[0] <= 1'b0;
                    stage2_col69[1] <= 1'b0;
                    stage2_col69[2] <= 1'b0;
                    stage2_col69[3] <= 1'b0;
                    stage2_col69[4] <= 1'b0;
                    stage2_col69[5] <= 1'b0;
                    stage2_col69[6] <= 1'b0;
                    stage2_col69[7] <= 1'b0;
                    stage2_col69[8] <= 1'b0;
                    stage2_col69[9] <= 1'b0;
                    stage2_col69[10] <= 1'b0;
                    stage2_col69[11] <= 1'b0;
                    stage2_col69[12] <= 1'b0;
                    stage2_col69[13] <= 1'b0;
                    stage2_col69[14] <= 1'b0;
                    stage2_col69[15] <= 1'b0;
                    stage2_col70[0] <= 1'b0;
                    stage2_col70[1] <= 1'b0;
                    stage2_col70[2] <= 1'b0;
                    stage2_col70[3] <= 1'b0;
                    stage2_col70[4] <= 1'b0;
                    stage2_col70[5] <= 1'b0;
                    stage2_col70[6] <= 1'b0;
                    stage2_col70[7] <= 1'b0;
                    stage2_col70[8] <= 1'b0;
                    stage2_col70[9] <= 1'b0;
                    stage2_col70[10] <= 1'b0;
                    stage2_col70[11] <= 1'b0;
                    stage2_col70[12] <= 1'b0;
                    stage2_col70[13] <= 1'b0;
                    stage2_col71[0] <= 1'b0;
                    stage2_col71[1] <= 1'b0;
                    stage2_col71[2] <= 1'b0;
                    stage2_col71[3] <= 1'b0;
                    stage2_col71[4] <= 1'b0;
                    stage2_col71[5] <= 1'b0;
                    stage2_col71[6] <= 1'b0;
                    stage2_col71[7] <= 1'b0;
                    stage2_col71[8] <= 1'b0;
                    stage2_col71[9] <= 1'b0;
                    stage2_col71[10] <= 1'b0;
                    stage2_col71[11] <= 1'b0;
                    stage2_col71[12] <= 1'b0;
                    stage2_col71[13] <= 1'b0;
                    stage2_col71[14] <= 1'b0;
                    stage2_col71[15] <= 1'b0;
                    stage2_col72[0] <= 1'b0;
                    stage2_col72[1] <= 1'b0;
                    stage2_col72[2] <= 1'b0;
                    stage2_col72[3] <= 1'b0;
                    stage2_col72[4] <= 1'b0;
                    stage2_col72[5] <= 1'b0;
                    stage2_col72[6] <= 1'b0;
                    stage2_col72[7] <= 1'b0;
                    stage2_col72[8] <= 1'b0;
                    stage2_col72[9] <= 1'b0;
                    stage2_col72[10] <= 1'b0;
                    stage2_col72[11] <= 1'b0;
                    stage2_col72[12] <= 1'b0;
                    stage2_col72[13] <= 1'b0;
                    stage2_col73[0] <= 1'b0;
                    stage2_col73[1] <= 1'b0;
                    stage2_col73[2] <= 1'b0;
                    stage2_col73[3] <= 1'b0;
                    stage2_col73[4] <= 1'b0;
                    stage2_col73[5] <= 1'b0;
                    stage2_col73[6] <= 1'b0;
                    stage2_col73[7] <= 1'b0;
                    stage2_col73[8] <= 1'b0;
                    stage2_col73[9] <= 1'b0;
                    stage2_col73[10] <= 1'b0;
                    stage2_col73[11] <= 1'b0;
                    stage2_col73[12] <= 1'b0;
                    stage2_col73[13] <= 1'b0;
                    stage2_col73[14] <= 1'b0;
                    stage2_col73[15] <= 1'b0;
                    stage2_col74[0] <= 1'b0;
                    stage2_col74[1] <= 1'b0;
                    stage2_col74[2] <= 1'b0;
                    stage2_col74[3] <= 1'b0;
                    stage2_col74[4] <= 1'b0;
                    stage2_col74[5] <= 1'b0;
                    stage2_col74[6] <= 1'b0;
                    stage2_col74[7] <= 1'b0;
                    stage2_col74[8] <= 1'b0;
                    stage2_col74[9] <= 1'b0;
                    stage2_col74[10] <= 1'b0;
                    stage2_col74[11] <= 1'b0;
                    stage2_col74[12] <= 1'b0;
                    stage2_col74[13] <= 1'b0;
                    stage2_col75[0] <= 1'b0;
                    stage2_col75[1] <= 1'b0;
                    stage2_col75[2] <= 1'b0;
                    stage2_col75[3] <= 1'b0;
                    stage2_col75[4] <= 1'b0;
                    stage2_col75[5] <= 1'b0;
                    stage2_col75[6] <= 1'b0;
                    stage2_col75[7] <= 1'b0;
                    stage2_col75[8] <= 1'b0;
                    stage2_col75[9] <= 1'b0;
                    stage2_col75[10] <= 1'b0;
                    stage2_col75[11] <= 1'b0;
                    stage2_col75[12] <= 1'b0;
                    stage2_col75[13] <= 1'b0;
                    stage2_col75[14] <= 1'b0;
                    stage2_col75[15] <= 1'b0;
                    stage2_col76[0] <= 1'b0;
                    stage2_col76[1] <= 1'b0;
                    stage2_col76[2] <= 1'b0;
                    stage2_col76[3] <= 1'b0;
                    stage2_col76[4] <= 1'b0;
                    stage2_col76[5] <= 1'b0;
                    stage2_col76[6] <= 1'b0;
                    stage2_col76[7] <= 1'b0;
                    stage2_col76[8] <= 1'b0;
                    stage2_col76[9] <= 1'b0;
                    stage2_col76[10] <= 1'b0;
                    stage2_col76[11] <= 1'b0;
                    stage2_col76[12] <= 1'b0;
                    stage2_col76[13] <= 1'b0;
                    stage2_col77[0] <= 1'b0;
                    stage2_col77[1] <= 1'b0;
                    stage2_col77[2] <= 1'b0;
                    stage2_col77[3] <= 1'b0;
                    stage2_col77[4] <= 1'b0;
                    stage2_col77[5] <= 1'b0;
                    stage2_col77[6] <= 1'b0;
                    stage2_col77[7] <= 1'b0;
                    stage2_col77[8] <= 1'b0;
                    stage2_col77[9] <= 1'b0;
                    stage2_col77[10] <= 1'b0;
                    stage2_col77[11] <= 1'b0;
                    stage2_col77[12] <= 1'b0;
                    stage2_col77[13] <= 1'b0;
                    stage2_col77[14] <= 1'b0;
                    stage2_col77[15] <= 1'b0;
                    stage2_col78[0] <= 1'b0;
                    stage2_col78[1] <= 1'b0;
                    stage2_col78[2] <= 1'b0;
                    stage2_col78[3] <= 1'b0;
                    stage2_col78[4] <= 1'b0;
                    stage2_col78[5] <= 1'b0;
                    stage2_col78[6] <= 1'b0;
                    stage2_col78[7] <= 1'b0;
                    stage2_col78[8] <= 1'b0;
                    stage2_col78[9] <= 1'b0;
                    stage2_col78[10] <= 1'b0;
                    stage2_col78[11] <= 1'b0;
                    stage2_col78[12] <= 1'b0;
                    stage2_col78[13] <= 1'b0;
                    stage2_col79[0] <= 1'b0;
                    stage2_col79[1] <= 1'b0;
                    stage2_col79[2] <= 1'b0;
                    stage2_col79[3] <= 1'b0;
                    stage2_col79[4] <= 1'b0;
                    stage2_col79[5] <= 1'b0;
                    stage2_col79[6] <= 1'b0;
                    stage2_col79[7] <= 1'b0;
                    stage2_col79[8] <= 1'b0;
                    stage2_col79[9] <= 1'b0;
                    stage2_col79[10] <= 1'b0;
                    stage2_col79[11] <= 1'b0;
                    stage2_col79[12] <= 1'b0;
                    stage2_col79[13] <= 1'b0;
                    stage2_col79[14] <= 1'b0;
                    stage2_col79[15] <= 1'b0;
                    stage2_col80[0] <= 1'b0;
                    stage2_col80[1] <= 1'b0;
                    stage2_col80[2] <= 1'b0;
                    stage2_col80[3] <= 1'b0;
                    stage2_col80[4] <= 1'b0;
                    stage2_col80[5] <= 1'b0;
                    stage2_col80[6] <= 1'b0;
                    stage2_col80[7] <= 1'b0;
                    stage2_col80[8] <= 1'b0;
                    stage2_col80[9] <= 1'b0;
                    stage2_col80[10] <= 1'b0;
                    stage2_col80[11] <= 1'b0;
                    stage2_col80[12] <= 1'b0;
                    stage2_col80[13] <= 1'b0;
                    stage2_col81[0] <= 1'b0;
                    stage2_col81[1] <= 1'b0;
                    stage2_col81[2] <= 1'b0;
                    stage2_col81[3] <= 1'b0;
                    stage2_col81[4] <= 1'b0;
                    stage2_col81[5] <= 1'b0;
                    stage2_col81[6] <= 1'b0;
                    stage2_col81[7] <= 1'b0;
                    stage2_col81[8] <= 1'b0;
                    stage2_col81[9] <= 1'b0;
                    stage2_col81[10] <= 1'b0;
                    stage2_col81[11] <= 1'b0;
                    stage2_col81[12] <= 1'b0;
                    stage2_col81[13] <= 1'b0;
                    stage2_col81[14] <= 1'b0;
                    stage2_col81[15] <= 1'b0;
                    stage2_col82[0] <= 1'b0;
                    stage2_col82[1] <= 1'b0;
                    stage2_col82[2] <= 1'b0;
                    stage2_col82[3] <= 1'b0;
                    stage2_col82[4] <= 1'b0;
                    stage2_col82[5] <= 1'b0;
                    stage2_col82[6] <= 1'b0;
                    stage2_col82[7] <= 1'b0;
                    stage2_col82[8] <= 1'b0;
                    stage2_col82[9] <= 1'b0;
                    stage2_col82[10] <= 1'b0;
                    stage2_col82[11] <= 1'b0;
                    stage2_col82[12] <= 1'b0;
                    stage2_col82[13] <= 1'b0;
                    stage2_col83[0] <= 1'b0;
                    stage2_col83[1] <= 1'b0;
                    stage2_col83[2] <= 1'b0;
                    stage2_col83[3] <= 1'b0;
                    stage2_col83[4] <= 1'b0;
                    stage2_col83[5] <= 1'b0;
                    stage2_col83[6] <= 1'b0;
                    stage2_col83[7] <= 1'b0;
                    stage2_col83[8] <= 1'b0;
                    stage2_col83[9] <= 1'b0;
                    stage2_col83[10] <= 1'b0;
                    stage2_col83[11] <= 1'b0;
                    stage2_col83[12] <= 1'b0;
                    stage2_col83[13] <= 1'b0;
                    stage2_col83[14] <= 1'b0;
                    stage2_col83[15] <= 1'b0;
                    stage2_col84[0] <= 1'b0;
                    stage2_col84[1] <= 1'b0;
                    stage2_col84[2] <= 1'b0;
                    stage2_col84[3] <= 1'b0;
                    stage2_col84[4] <= 1'b0;
                    stage2_col84[5] <= 1'b0;
                    stage2_col84[6] <= 1'b0;
                    stage2_col84[7] <= 1'b0;
                    stage2_col84[8] <= 1'b0;
                    stage2_col84[9] <= 1'b0;
                    stage2_col84[10] <= 1'b0;
                    stage2_col84[11] <= 1'b0;
                    stage2_col84[12] <= 1'b0;
                    stage2_col84[13] <= 1'b0;
                    stage2_col85[0] <= 1'b0;
                    stage2_col85[1] <= 1'b0;
                    stage2_col85[2] <= 1'b0;
                    stage2_col85[3] <= 1'b0;
                    stage2_col85[4] <= 1'b0;
                    stage2_col85[5] <= 1'b0;
                    stage2_col85[6] <= 1'b0;
                    stage2_col85[7] <= 1'b0;
                    stage2_col85[8] <= 1'b0;
                    stage2_col85[9] <= 1'b0;
                    stage2_col85[10] <= 1'b0;
                    stage2_col85[11] <= 1'b0;
                    stage2_col85[12] <= 1'b0;
                    stage2_col85[13] <= 1'b0;
                    stage2_col85[14] <= 1'b0;
                    stage2_col85[15] <= 1'b0;
                    stage2_col86[0] <= 1'b0;
                    stage2_col86[1] <= 1'b0;
                    stage2_col86[2] <= 1'b0;
                    stage2_col86[3] <= 1'b0;
                    stage2_col86[4] <= 1'b0;
                    stage2_col86[5] <= 1'b0;
                    stage2_col86[6] <= 1'b0;
                    stage2_col86[7] <= 1'b0;
                    stage2_col86[8] <= 1'b0;
                    stage2_col86[9] <= 1'b0;
                    stage2_col86[10] <= 1'b0;
                    stage2_col86[11] <= 1'b0;
                    stage2_col86[12] <= 1'b0;
                    stage2_col86[13] <= 1'b0;
                    stage2_col87[0] <= 1'b0;
                    stage2_col87[1] <= 1'b0;
                    stage2_col87[2] <= 1'b0;
                    stage2_col87[3] <= 1'b0;
                    stage2_col87[4] <= 1'b0;
                    stage2_col87[5] <= 1'b0;
                    stage2_col87[6] <= 1'b0;
                    stage2_col87[7] <= 1'b0;
                    stage2_col87[8] <= 1'b0;
                    stage2_col87[9] <= 1'b0;
                    stage2_col87[10] <= 1'b0;
                    stage2_col87[11] <= 1'b0;
                    stage2_col87[12] <= 1'b0;
                    stage2_col87[13] <= 1'b0;
                    stage2_col87[14] <= 1'b0;
                    stage2_col87[15] <= 1'b0;
                    stage2_col88[0] <= 1'b0;
                    stage2_col88[1] <= 1'b0;
                    stage2_col88[2] <= 1'b0;
                    stage2_col88[3] <= 1'b0;
                    stage2_col88[4] <= 1'b0;
                    stage2_col88[5] <= 1'b0;
                    stage2_col88[6] <= 1'b0;
                    stage2_col88[7] <= 1'b0;
                    stage2_col88[8] <= 1'b0;
                    stage2_col88[9] <= 1'b0;
                    stage2_col88[10] <= 1'b0;
                    stage2_col88[11] <= 1'b0;
                    stage2_col88[12] <= 1'b0;
                    stage2_col88[13] <= 1'b0;
                    stage2_col89[0] <= 1'b0;
                    stage2_col89[1] <= 1'b0;
                    stage2_col89[2] <= 1'b0;
                    stage2_col89[3] <= 1'b0;
                    stage2_col89[4] <= 1'b0;
                    stage2_col89[5] <= 1'b0;
                    stage2_col89[6] <= 1'b0;
                    stage2_col89[7] <= 1'b0;
                    stage2_col89[8] <= 1'b0;
                    stage2_col89[9] <= 1'b0;
                    stage2_col89[10] <= 1'b0;
                    stage2_col89[11] <= 1'b0;
                    stage2_col89[12] <= 1'b0;
                    stage2_col89[13] <= 1'b0;
                    stage2_col89[14] <= 1'b0;
                    stage2_col89[15] <= 1'b0;
                    stage2_col90[0] <= 1'b0;
                    stage2_col90[1] <= 1'b0;
                    stage2_col90[2] <= 1'b0;
                    stage2_col90[3] <= 1'b0;
                    stage2_col90[4] <= 1'b0;
                    stage2_col90[5] <= 1'b0;
                    stage2_col90[6] <= 1'b0;
                    stage2_col90[7] <= 1'b0;
                    stage2_col90[8] <= 1'b0;
                    stage2_col90[9] <= 1'b0;
                    stage2_col90[10] <= 1'b0;
                    stage2_col90[11] <= 1'b0;
                    stage2_col90[12] <= 1'b0;
                    stage2_col90[13] <= 1'b0;
                    stage2_col91[0] <= 1'b0;
                    stage2_col91[1] <= 1'b0;
                    stage2_col91[2] <= 1'b0;
                    stage2_col91[3] <= 1'b0;
                    stage2_col91[4] <= 1'b0;
                    stage2_col91[5] <= 1'b0;
                    stage2_col91[6] <= 1'b0;
                    stage2_col91[7] <= 1'b0;
                    stage2_col91[8] <= 1'b0;
                    stage2_col91[9] <= 1'b0;
                    stage2_col91[10] <= 1'b0;
                    stage2_col91[11] <= 1'b0;
                    stage2_col91[12] <= 1'b0;
                    stage2_col91[13] <= 1'b0;
                    stage2_col91[14] <= 1'b0;
                    stage2_col91[15] <= 1'b0;
                    stage2_col92[0] <= 1'b0;
                    stage2_col92[1] <= 1'b0;
                    stage2_col92[2] <= 1'b0;
                    stage2_col92[3] <= 1'b0;
                    stage2_col92[4] <= 1'b0;
                    stage2_col92[5] <= 1'b0;
                    stage2_col92[6] <= 1'b0;
                    stage2_col92[7] <= 1'b0;
                    stage2_col92[8] <= 1'b0;
                    stage2_col92[9] <= 1'b0;
                    stage2_col92[10] <= 1'b0;
                    stage2_col92[11] <= 1'b0;
                    stage2_col92[12] <= 1'b0;
                    stage2_col92[13] <= 1'b0;
                    stage2_col93[0] <= 1'b0;
                    stage2_col93[1] <= 1'b0;
                    stage2_col93[2] <= 1'b0;
                    stage2_col93[3] <= 1'b0;
                    stage2_col93[4] <= 1'b0;
                    stage2_col93[5] <= 1'b0;
                    stage2_col93[6] <= 1'b0;
                    stage2_col93[7] <= 1'b0;
                    stage2_col93[8] <= 1'b0;
                    stage2_col93[9] <= 1'b0;
                    stage2_col93[10] <= 1'b0;
                    stage2_col93[11] <= 1'b0;
                    stage2_col93[12] <= 1'b0;
                    stage2_col93[13] <= 1'b0;
                    stage2_col93[14] <= 1'b0;
                    stage2_col93[15] <= 1'b0;
                    stage2_col94[0] <= 1'b0;
                    stage2_col94[1] <= 1'b0;
                    stage2_col94[2] <= 1'b0;
                    stage2_col94[3] <= 1'b0;
                    stage2_col94[4] <= 1'b0;
                    stage2_col94[5] <= 1'b0;
                    stage2_col94[6] <= 1'b0;
                    stage2_col94[7] <= 1'b0;
                    stage2_col94[8] <= 1'b0;
                    stage2_col94[9] <= 1'b0;
                    stage2_col94[10] <= 1'b0;
                    stage2_col94[11] <= 1'b0;
                    stage2_col94[12] <= 1'b0;
                    stage2_col94[13] <= 1'b0;
                    stage2_col95[0] <= 1'b0;
                    stage2_col95[1] <= 1'b0;
                    stage2_col95[2] <= 1'b0;
                    stage2_col95[3] <= 1'b0;
                    stage2_col95[4] <= 1'b0;
                    stage2_col95[5] <= 1'b0;
                    stage2_col95[6] <= 1'b0;
                    stage2_col95[7] <= 1'b0;
                    stage2_col95[8] <= 1'b0;
                    stage2_col95[9] <= 1'b0;
                    stage2_col95[10] <= 1'b0;
                    stage2_col95[11] <= 1'b0;
                    stage2_col95[12] <= 1'b0;
                    stage2_col95[13] <= 1'b0;
                    stage2_col95[14] <= 1'b0;
                    stage2_col95[15] <= 1'b0;
                    stage2_col96[0] <= 1'b0;
                    stage2_col96[1] <= 1'b0;
                    stage2_col96[2] <= 1'b0;
                    stage2_col96[3] <= 1'b0;
                    stage2_col96[4] <= 1'b0;
                    stage2_col96[5] <= 1'b0;
                    stage2_col96[6] <= 1'b0;
                    stage2_col96[7] <= 1'b0;
                    stage2_col96[8] <= 1'b0;
                    stage2_col96[9] <= 1'b0;
                    stage2_col96[10] <= 1'b0;
                    stage2_col96[11] <= 1'b0;
                    stage2_col96[12] <= 1'b0;
                    stage2_col96[13] <= 1'b0;
                    stage2_col97[0] <= 1'b0;
                    stage2_col97[1] <= 1'b0;
                    stage2_col97[2] <= 1'b0;
                    stage2_col97[3] <= 1'b0;
                    stage2_col97[4] <= 1'b0;
                    stage2_col97[5] <= 1'b0;
                    stage2_col97[6] <= 1'b0;
                    stage2_col97[7] <= 1'b0;
                    stage2_col97[8] <= 1'b0;
                    stage2_col97[9] <= 1'b0;
                    stage2_col97[10] <= 1'b0;
                    stage2_col97[11] <= 1'b0;
                    stage2_col97[12] <= 1'b0;
                    stage2_col97[13] <= 1'b0;
                    stage2_col97[14] <= 1'b0;
                    stage2_col97[15] <= 1'b0;
                    stage2_col98[0] <= 1'b0;
                    stage2_col98[1] <= 1'b0;
                    stage2_col98[2] <= 1'b0;
                    stage2_col98[3] <= 1'b0;
                    stage2_col98[4] <= 1'b0;
                    stage2_col98[5] <= 1'b0;
                    stage2_col98[6] <= 1'b0;
                    stage2_col98[7] <= 1'b0;
                    stage2_col98[8] <= 1'b0;
                    stage2_col98[9] <= 1'b0;
                    stage2_col98[10] <= 1'b0;
                    stage2_col98[11] <= 1'b0;
                    stage2_col98[12] <= 1'b0;
                    stage2_col98[13] <= 1'b0;
                    stage2_col99[0] <= 1'b0;
                    stage2_col99[1] <= 1'b0;
                    stage2_col99[2] <= 1'b0;
                    stage2_col99[3] <= 1'b0;
                    stage2_col99[4] <= 1'b0;
                    stage2_col99[5] <= 1'b0;
                    stage2_col99[6] <= 1'b0;
                    stage2_col99[7] <= 1'b0;
                    stage2_col99[8] <= 1'b0;
                    stage2_col99[9] <= 1'b0;
                    stage2_col99[10] <= 1'b0;
                    stage2_col99[11] <= 1'b0;
                    stage2_col99[12] <= 1'b0;
                    stage2_col99[13] <= 1'b0;
                    stage2_col99[14] <= 1'b0;
                    stage2_col99[15] <= 1'b0;
                    stage2_col100[0] <= 1'b0;
                    stage2_col100[1] <= 1'b0;
                    stage2_col100[2] <= 1'b0;
                    stage2_col100[3] <= 1'b0;
                    stage2_col100[4] <= 1'b0;
                    stage2_col100[5] <= 1'b0;
                    stage2_col100[6] <= 1'b0;
                    stage2_col100[7] <= 1'b0;
                    stage2_col100[8] <= 1'b0;
                    stage2_col100[9] <= 1'b0;
                    stage2_col100[10] <= 1'b0;
                    stage2_col100[11] <= 1'b0;
                    stage2_col100[12] <= 1'b0;
                    stage2_col100[13] <= 1'b0;
                    stage2_col101[0] <= 1'b0;
                    stage2_col101[1] <= 1'b0;
                    stage2_col101[2] <= 1'b0;
                    stage2_col101[3] <= 1'b0;
                    stage2_col101[4] <= 1'b0;
                    stage2_col101[5] <= 1'b0;
                    stage2_col101[6] <= 1'b0;
                    stage2_col101[7] <= 1'b0;
                    stage2_col101[8] <= 1'b0;
                    stage2_col101[9] <= 1'b0;
                    stage2_col101[10] <= 1'b0;
                    stage2_col101[11] <= 1'b0;
                    stage2_col101[12] <= 1'b0;
                    stage2_col101[13] <= 1'b0;
                    stage2_col101[14] <= 1'b0;
                    stage2_col101[15] <= 1'b0;
                    stage2_col102[0] <= 1'b0;
                    stage2_col102[1] <= 1'b0;
                    stage2_col102[2] <= 1'b0;
                    stage2_col102[3] <= 1'b0;
                    stage2_col102[4] <= 1'b0;
                    stage2_col102[5] <= 1'b0;
                    stage2_col102[6] <= 1'b0;
                    stage2_col102[7] <= 1'b0;
                    stage2_col102[8] <= 1'b0;
                    stage2_col102[9] <= 1'b0;
                    stage2_col102[10] <= 1'b0;
                    stage2_col102[11] <= 1'b0;
                    stage2_col102[12] <= 1'b0;
                    stage2_col102[13] <= 1'b0;
                    stage2_col103[0] <= 1'b0;
                    stage2_col103[1] <= 1'b0;
                    stage2_col103[2] <= 1'b0;
                    stage2_col103[3] <= 1'b0;
                    stage2_col103[4] <= 1'b0;
                    stage2_col103[5] <= 1'b0;
                    stage2_col103[6] <= 1'b0;
                    stage2_col103[7] <= 1'b0;
                    stage2_col103[8] <= 1'b0;
                    stage2_col103[9] <= 1'b0;
                    stage2_col103[10] <= 1'b0;
                    stage2_col103[11] <= 1'b0;
                    stage2_col103[12] <= 1'b0;
                    stage2_col103[13] <= 1'b0;
                    stage2_col103[14] <= 1'b0;
                    stage2_col103[15] <= 1'b0;
                    stage2_col104[0] <= 1'b0;
                    stage2_col104[1] <= 1'b0;
                    stage2_col104[2] <= 1'b0;
                    stage2_col104[3] <= 1'b0;
                    stage2_col104[4] <= 1'b0;
                    stage2_col104[5] <= 1'b0;
                    stage2_col104[6] <= 1'b0;
                    stage2_col104[7] <= 1'b0;
                    stage2_col104[8] <= 1'b0;
                    stage2_col104[9] <= 1'b0;
                    stage2_col104[10] <= 1'b0;
                    stage2_col104[11] <= 1'b0;
                    stage2_col104[12] <= 1'b0;
                    stage2_col104[13] <= 1'b0;
                    stage2_col105[0] <= 1'b0;
                    stage2_col105[1] <= 1'b0;
                    stage2_col105[2] <= 1'b0;
                    stage2_col105[3] <= 1'b0;
                    stage2_col105[4] <= 1'b0;
                    stage2_col105[5] <= 1'b0;
                    stage2_col105[6] <= 1'b0;
                    stage2_col105[7] <= 1'b0;
                    stage2_col105[8] <= 1'b0;
                    stage2_col105[9] <= 1'b0;
                    stage2_col105[10] <= 1'b0;
                    stage2_col105[11] <= 1'b0;
                    stage2_col105[12] <= 1'b0;
                    stage2_col105[13] <= 1'b0;
                    stage2_col105[14] <= 1'b0;
                    stage2_col105[15] <= 1'b0;
                    stage2_col106[0] <= 1'b0;
                    stage2_col106[1] <= 1'b0;
                    stage2_col106[2] <= 1'b0;
                    stage2_col106[3] <= 1'b0;
                    stage2_col106[4] <= 1'b0;
                    stage2_col106[5] <= 1'b0;
                    stage2_col106[6] <= 1'b0;
                    stage2_col106[7] <= 1'b0;
                    stage2_col106[8] <= 1'b0;
                    stage2_col106[9] <= 1'b0;
                    stage2_col106[10] <= 1'b0;
                    stage2_col106[11] <= 1'b0;
                    stage2_col106[12] <= 1'b0;
                    stage2_col106[13] <= 1'b0;
                    stage2_col107[0] <= 1'b0;
                    stage2_col107[1] <= 1'b0;
                    stage2_col107[2] <= 1'b0;
                    stage2_col107[3] <= 1'b0;
                    stage2_col107[4] <= 1'b0;
                    stage2_col107[5] <= 1'b0;
                    stage2_col107[6] <= 1'b0;
                    stage2_col107[7] <= 1'b0;
                    stage2_col107[8] <= 1'b0;
                    stage2_col107[9] <= 1'b0;
                    stage2_col107[10] <= 1'b0;
                    stage2_col107[11] <= 1'b0;
                    stage2_col107[12] <= 1'b0;
                    stage2_col107[13] <= 1'b0;
                    stage2_col107[14] <= 1'b0;
                    stage2_col107[15] <= 1'b0;
                    stage2_col108[0] <= 1'b0;
                    stage2_col108[1] <= 1'b0;
                    stage2_col108[2] <= 1'b0;
                    stage2_col108[3] <= 1'b0;
                    stage2_col108[4] <= 1'b0;
                    stage2_col108[5] <= 1'b0;
                    stage2_col108[6] <= 1'b0;
                    stage2_col108[7] <= 1'b0;
                    stage2_col108[8] <= 1'b0;
                    stage2_col108[9] <= 1'b0;
                    stage2_col108[10] <= 1'b0;
                    stage2_col108[11] <= 1'b0;
                    stage2_col108[12] <= 1'b0;
                    stage2_col108[13] <= 1'b0;
                    stage2_col109[0] <= 1'b0;
                    stage2_col109[1] <= 1'b0;
                    stage2_col109[2] <= 1'b0;
                    stage2_col109[3] <= 1'b0;
                    stage2_col109[4] <= 1'b0;
                    stage2_col109[5] <= 1'b0;
                    stage2_col109[6] <= 1'b0;
                    stage2_col109[7] <= 1'b0;
                    stage2_col109[8] <= 1'b0;
                    stage2_col109[9] <= 1'b0;
                    stage2_col109[10] <= 1'b0;
                    stage2_col109[11] <= 1'b0;
                    stage2_col109[12] <= 1'b0;
                    stage2_col109[13] <= 1'b0;
                    stage2_col109[14] <= 1'b0;
                    stage2_col109[15] <= 1'b0;
                    stage2_col110[0] <= 1'b0;
                    stage2_col110[1] <= 1'b0;
                    stage2_col110[2] <= 1'b0;
                    stage2_col110[3] <= 1'b0;
                    stage2_col110[4] <= 1'b0;
                    stage2_col110[5] <= 1'b0;
                    stage2_col110[6] <= 1'b0;
                    stage2_col110[7] <= 1'b0;
                    stage2_col110[8] <= 1'b0;
                    stage2_col110[9] <= 1'b0;
                    stage2_col110[10] <= 1'b0;
                    stage2_col110[11] <= 1'b0;
                    stage2_col110[12] <= 1'b0;
                    stage2_col110[13] <= 1'b0;
                    stage2_col111[0] <= 1'b0;
                    stage2_col111[1] <= 1'b0;
                    stage2_col111[2] <= 1'b0;
                    stage2_col111[3] <= 1'b0;
                    stage2_col111[4] <= 1'b0;
                    stage2_col111[5] <= 1'b0;
                    stage2_col111[6] <= 1'b0;
                    stage2_col111[7] <= 1'b0;
                    stage2_col111[8] <= 1'b0;
                    stage2_col111[9] <= 1'b0;
                    stage2_col111[10] <= 1'b0;
                    stage2_col111[11] <= 1'b0;
                    stage2_col111[12] <= 1'b0;
                    stage2_col111[13] <= 1'b0;
                    stage2_col111[14] <= 1'b0;
                    stage2_col111[15] <= 1'b0;
                    stage2_col112[0] <= 1'b0;
                    stage2_col112[1] <= 1'b0;
                    stage2_col112[2] <= 1'b0;
                    stage2_col112[3] <= 1'b0;
                    stage2_col112[4] <= 1'b0;
                    stage2_col112[5] <= 1'b0;
                    stage2_col112[6] <= 1'b0;
                    stage2_col112[7] <= 1'b0;
                    stage2_col112[8] <= 1'b0;
                    stage2_col112[9] <= 1'b0;
                    stage2_col112[10] <= 1'b0;
                    stage2_col112[11] <= 1'b0;
                    stage2_col112[12] <= 1'b0;
                    stage2_col112[13] <= 1'b0;
                    stage2_col113[0] <= 1'b0;
                    stage2_col113[1] <= 1'b0;
                    stage2_col113[2] <= 1'b0;
                    stage2_col113[3] <= 1'b0;
                    stage2_col113[4] <= 1'b0;
                    stage2_col113[5] <= 1'b0;
                    stage2_col113[6] <= 1'b0;
                    stage2_col113[7] <= 1'b0;
                    stage2_col113[8] <= 1'b0;
                    stage2_col113[9] <= 1'b0;
                    stage2_col113[10] <= 1'b0;
                    stage2_col113[11] <= 1'b0;
                    stage2_col113[12] <= 1'b0;
                    stage2_col113[13] <= 1'b0;
                    stage2_col113[14] <= 1'b0;
                    stage2_col113[15] <= 1'b0;
                    stage2_col114[0] <= 1'b0;
                    stage2_col114[1] <= 1'b0;
                    stage2_col114[2] <= 1'b0;
                    stage2_col114[3] <= 1'b0;
                    stage2_col114[4] <= 1'b0;
                    stage2_col114[5] <= 1'b0;
                    stage2_col114[6] <= 1'b0;
                    stage2_col114[7] <= 1'b0;
                    stage2_col114[8] <= 1'b0;
                    stage2_col114[9] <= 1'b0;
                    stage2_col114[10] <= 1'b0;
                    stage2_col114[11] <= 1'b0;
                    stage2_col114[12] <= 1'b0;
                    stage2_col114[13] <= 1'b0;
                    stage2_col115[0] <= 1'b0;
                    stage2_col115[1] <= 1'b0;
                    stage2_col115[2] <= 1'b0;
                    stage2_col115[3] <= 1'b0;
                    stage2_col115[4] <= 1'b0;
                    stage2_col115[5] <= 1'b0;
                    stage2_col115[6] <= 1'b0;
                    stage2_col115[7] <= 1'b0;
                    stage2_col115[8] <= 1'b0;
                    stage2_col115[9] <= 1'b0;
                    stage2_col115[10] <= 1'b0;
                    stage2_col115[11] <= 1'b0;
                    stage2_col115[12] <= 1'b0;
                    stage2_col115[13] <= 1'b0;
                    stage2_col115[14] <= 1'b0;
                    stage2_col115[15] <= 1'b0;
                    stage2_col116[0] <= 1'b0;
                    stage2_col116[1] <= 1'b0;
                    stage2_col116[2] <= 1'b0;
                    stage2_col116[3] <= 1'b0;
                    stage2_col116[4] <= 1'b0;
                    stage2_col116[5] <= 1'b0;
                    stage2_col116[6] <= 1'b0;
                    stage2_col116[7] <= 1'b0;
                    stage2_col116[8] <= 1'b0;
                    stage2_col116[9] <= 1'b0;
                    stage2_col116[10] <= 1'b0;
                    stage2_col116[11] <= 1'b0;
                    stage2_col116[12] <= 1'b0;
                    stage2_col116[13] <= 1'b0;
                    stage2_col117[0] <= 1'b0;
                    stage2_col117[1] <= 1'b0;
                    stage2_col117[2] <= 1'b0;
                    stage2_col117[3] <= 1'b0;
                    stage2_col117[4] <= 1'b0;
                    stage2_col117[5] <= 1'b0;
                    stage2_col117[6] <= 1'b0;
                    stage2_col117[7] <= 1'b0;
                    stage2_col117[8] <= 1'b0;
                    stage2_col117[9] <= 1'b0;
                    stage2_col117[10] <= 1'b0;
                    stage2_col117[11] <= 1'b0;
                    stage2_col117[12] <= 1'b0;
                    stage2_col117[13] <= 1'b0;
                    stage2_col117[14] <= 1'b0;
                    stage2_col117[15] <= 1'b0;
                    stage2_col118[0] <= 1'b0;
                    stage2_col118[1] <= 1'b0;
                    stage2_col118[2] <= 1'b0;
                    stage2_col118[3] <= 1'b0;
                    stage2_col118[4] <= 1'b0;
                    stage2_col118[5] <= 1'b0;
                    stage2_col118[6] <= 1'b0;
                    stage2_col118[7] <= 1'b0;
                    stage2_col118[8] <= 1'b0;
                    stage2_col118[9] <= 1'b0;
                    stage2_col118[10] <= 1'b0;
                    stage2_col118[11] <= 1'b0;
                    stage2_col118[12] <= 1'b0;
                    stage2_col118[13] <= 1'b0;
                    stage2_col119[0] <= 1'b0;
                    stage2_col119[1] <= 1'b0;
                    stage2_col119[2] <= 1'b0;
                    stage2_col119[3] <= 1'b0;
                    stage2_col119[4] <= 1'b0;
                    stage2_col119[5] <= 1'b0;
                    stage2_col119[6] <= 1'b0;
                    stage2_col119[7] <= 1'b0;
                    stage2_col119[8] <= 1'b0;
                    stage2_col119[9] <= 1'b0;
                    stage2_col119[10] <= 1'b0;
                    stage2_col119[11] <= 1'b0;
                    stage2_col119[12] <= 1'b0;
                    stage2_col119[13] <= 1'b0;
                    stage2_col119[14] <= 1'b0;
                    stage2_col119[15] <= 1'b0;
                    stage2_col120[0] <= 1'b0;
                    stage2_col120[1] <= 1'b0;
                    stage2_col120[2] <= 1'b0;
                    stage2_col120[3] <= 1'b0;
                    stage2_col120[4] <= 1'b0;
                    stage2_col120[5] <= 1'b0;
                    stage2_col120[6] <= 1'b0;
                    stage2_col120[7] <= 1'b0;
                    stage2_col120[8] <= 1'b0;
                    stage2_col120[9] <= 1'b0;
                    stage2_col120[10] <= 1'b0;
                    stage2_col120[11] <= 1'b0;
                    stage2_col120[12] <= 1'b0;
                    stage2_col120[13] <= 1'b0;
                    stage2_col121[0] <= 1'b0;
                    stage2_col121[1] <= 1'b0;
                    stage2_col121[2] <= 1'b0;
                    stage2_col121[3] <= 1'b0;
                    stage2_col121[4] <= 1'b0;
                    stage2_col121[5] <= 1'b0;
                    stage2_col121[6] <= 1'b0;
                    stage2_col121[7] <= 1'b0;
                    stage2_col121[8] <= 1'b0;
                    stage2_col121[9] <= 1'b0;
                    stage2_col121[10] <= 1'b0;
                    stage2_col121[11] <= 1'b0;
                    stage2_col121[12] <= 1'b0;
                    stage2_col121[13] <= 1'b0;
                    stage2_col121[14] <= 1'b0;
                    stage2_col121[15] <= 1'b0;
                    stage2_col122[0] <= 1'b0;
                    stage2_col122[1] <= 1'b0;
                    stage2_col122[2] <= 1'b0;
                    stage2_col122[3] <= 1'b0;
                    stage2_col122[4] <= 1'b0;
                    stage2_col122[5] <= 1'b0;
                    stage2_col122[6] <= 1'b0;
                    stage2_col122[7] <= 1'b0;
                    stage2_col122[8] <= 1'b0;
                    stage2_col122[9] <= 1'b0;
                    stage2_col122[10] <= 1'b0;
                    stage2_col122[11] <= 1'b0;
                    stage2_col122[12] <= 1'b0;
                    stage2_col122[13] <= 1'b0;
                    stage2_col123[0] <= 1'b0;
                    stage2_col123[1] <= 1'b0;
                    stage2_col123[2] <= 1'b0;
                    stage2_col123[3] <= 1'b0;
                    stage2_col123[4] <= 1'b0;
                    stage2_col123[5] <= 1'b0;
                    stage2_col123[6] <= 1'b0;
                    stage2_col123[7] <= 1'b0;
                    stage2_col123[8] <= 1'b0;
                    stage2_col123[9] <= 1'b0;
                    stage2_col123[10] <= 1'b0;
                    stage2_col123[11] <= 1'b0;
                    stage2_col123[12] <= 1'b0;
                    stage2_col123[13] <= 1'b0;
                    stage2_col123[14] <= 1'b0;
                    stage2_col123[15] <= 1'b0;
                    stage2_col124[0] <= 1'b0;
                    stage2_col124[1] <= 1'b0;
                    stage2_col124[2] <= 1'b0;
                    stage2_col124[3] <= 1'b0;
                    stage2_col124[4] <= 1'b0;
                    stage2_col124[5] <= 1'b0;
                    stage2_col124[6] <= 1'b0;
                    stage2_col124[7] <= 1'b0;
                    stage2_col124[8] <= 1'b0;
                    stage2_col124[9] <= 1'b0;
                    stage2_col124[10] <= 1'b0;
                    stage2_col124[11] <= 1'b0;
                    stage2_col124[12] <= 1'b0;
                    stage2_col124[13] <= 1'b0;
                    stage2_col125[0] <= 1'b0;
                    stage2_col125[1] <= 1'b0;
                    stage2_col125[2] <= 1'b0;
                    stage2_col125[3] <= 1'b0;
                    stage2_col125[4] <= 1'b0;
                    stage2_col125[5] <= 1'b0;
                    stage2_col125[6] <= 1'b0;
                    stage2_col125[7] <= 1'b0;
                    stage2_col125[8] <= 1'b0;
                    stage2_col125[9] <= 1'b0;
                    stage2_col125[10] <= 1'b0;
                    stage2_col125[11] <= 1'b0;
                    stage2_col125[12] <= 1'b0;
                    stage2_col125[13] <= 1'b0;
                    stage2_col125[14] <= 1'b0;
                    stage2_col125[15] <= 1'b0;
                    stage2_col126[0] <= 1'b0;
                    stage2_col126[1] <= 1'b0;
                    stage2_col126[2] <= 1'b0;
                    stage2_col126[3] <= 1'b0;
                    stage2_col126[4] <= 1'b0;
                    stage2_col126[5] <= 1'b0;
                    stage2_col126[6] <= 1'b0;
                    stage2_col126[7] <= 1'b0;
                    stage2_col126[8] <= 1'b0;
                    stage2_col126[9] <= 1'b0;
                    stage2_col126[10] <= 1'b0;
                    stage2_col126[11] <= 1'b0;
                    stage2_col126[12] <= 1'b0;
                    stage2_col126[13] <= 1'b0;
                    stage2_col127[0] <= 1'b0;
                    stage2_col127[1] <= 1'b0;
                    stage2_col127[2] <= 1'b0;
                    stage2_col127[3] <= 1'b0;
                    stage2_col127[4] <= 1'b0;
                    stage2_col127[5] <= 1'b0;
                    stage2_col127[6] <= 1'b0;
                    stage2_col127[7] <= 1'b0;
                    stage2_col127[8] <= 1'b0;
                    stage2_col127[9] <= 1'b0;
                    stage2_col127[10] <= 1'b0;
                    stage2_col127[11] <= 1'b0;
                    stage2_col127[12] <= 1'b0;
                    stage2_col127[13] <= 1'b0;
                    stage2_col127[14] <= 1'b0;
                    stage2_col127[15] <= 1'b0;
                    stage2_col127[16] <= 1'b0;
                    stage2_col127[17] <= 1'b0;
                    stage2_col127[18] <= 1'b0;
                    stage2_col127[19] <= 1'b0;
                    stage2_col127[20] <= 1'b0;
                    stage2_col127[21] <= 1'b0;
                    stage2_col127[22] <= 1'b0;
                    stage2_col127[23] <= 1'b0;
                    stage2_col127[24] <= 1'b0;
                    stage2_col127[25] <= 1'b0;
                    stage2_col127[26] <= 1'b0;
                    stage2_col127[27] <= 1'b0;
                    stage2_col127[28] <= 1'b0;
                    stage2_col127[29] <= 1'b0;
                    stage2_col127[30] <= 1'b0;
                    stage2_col127[31] <= 1'b0;
                    stage2_col127[32] <= 1'b0;
                    stage2_col127[33] <= 1'b0;
                    stage2_col127[34] <= 1'b0;
                    stage2_col127[35] <= 1'b0;
                    stage2_col127[36] <= 1'b0;
                    stage2_col127[37] <= 1'b0;
                    stage2_col127[38] <= 1'b0;
                    stage2_col127[39] <= 1'b0;
                    stage2_col127[40] <= 1'b0;
                    stage2_col127[41] <= 1'b0;
                    stage2_col127[42] <= 1'b0;
                    stage2_col127[43] <= 1'b0;
                    stage2_col127[44] <= 1'b0;
                    stage2_col127[45] <= 1'b0;
                    stage2_col127[46] <= 1'b0;
                    stage2_col127[47] <= 1'b0;
                    stage2_col127[48] <= 1'b0;
                    stage2_col127[49] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage2_col0[0] <= stage1_col0[0];
                    stage2_col1[0] <= ha_s1_c1_n0_s;
                    stage2_col2[0] <= ha_s1_c1_n0_c;
                    stage2_col2[1] <= stage1_col2[0];
                    stage2_col3[0] <= fa_s1_c3_n0_s;
                    stage2_col4[0] <= fa_s1_c3_n0_c;
                    stage2_col4[1] <= stage1_col4[0];
                    stage2_col4[2] <= stage1_col4[1];
                    stage2_col5[0] <= stage1_col5[0];
                    stage2_col5[1] <= stage1_col5[1];
                    stage2_col6[0] <= fa_s1_c6_n1_s;
                    stage2_col6[1] <= stage1_col6[3];
                    stage2_col7[0] <= fa_s1_c6_n1_c;
                    stage2_col7[1] <= fa_s1_c7_n2_s;
                    stage2_col8[0] <= fa_s1_c7_n2_c;
                    stage2_col8[1] <= fa_s1_c8_n3_s;
                    stage2_col9[0] <= fa_s1_c8_n3_c;
                    stage2_col9[1] <= fa_s1_c9_n4_s;
                    stage2_col9[2] <= stage1_col9[3];
                    stage2_col9[3] <= stage1_col9[4];
                    stage2_col10[0] <= fa_s1_c9_n4_c;
                    stage2_col10[1] <= fa_s1_c10_n5_s;
                    stage2_col10[2] <= stage1_col10[3];
                    stage2_col11[0] <= fa_s1_c10_n5_c;
                    stage2_col11[1] <= fa_s1_c11_n6_s;
                    stage2_col11[2] <= stage1_col11[3];
                    stage2_col12[0] <= fa_s1_c11_n6_c;
                    stage2_col12[1] <= fa_s1_c12_n7_s;
                    stage2_col12[2] <= fa_s1_c12_n8_s;
                    stage2_col13[0] <= fa_s1_c12_n7_c;
                    stage2_col13[1] <= fa_s1_c12_n8_c;
                    stage2_col13[2] <= fa_s1_c13_n9_s;
                    stage2_col13[3] <= stage1_col13[3];
                    stage2_col13[4] <= stage1_col13[4];
                    stage2_col14[0] <= fa_s1_c13_n9_c;
                    stage2_col14[1] <= fa_s1_c14_n10_s;
                    stage2_col14[2] <= stage1_col14[3];
                    stage2_col14[3] <= stage1_col14[4];
                    stage2_col15[0] <= fa_s1_c14_n10_c;
                    stage2_col15[1] <= fa_s1_c15_n11_s;
                    stage2_col15[2] <= fa_s1_c15_n12_s;
                    stage2_col15[3] <= stage1_col15[6];
                    stage2_col16[0] <= fa_s1_c15_n11_c;
                    stage2_col16[1] <= fa_s1_c15_n12_c;
                    stage2_col16[2] <= fa_s1_c16_n13_s;
                    stage2_col16[3] <= fa_s1_c16_n14_s;
                    stage2_col17[0] <= fa_s1_c16_n13_c;
                    stage2_col17[1] <= fa_s1_c16_n14_c;
                    stage2_col17[2] <= fa_s1_c17_n15_s;
                    stage2_col17[3] <= fa_s1_c17_n16_s;
                    stage2_col18[0] <= fa_s1_c17_n15_c;
                    stage2_col18[1] <= fa_s1_c17_n16_c;
                    stage2_col18[2] <= fa_s1_c18_n17_s;
                    stage2_col18[3] <= fa_s1_c18_n18_s;
                    stage2_col18[4] <= stage1_col18[6];
                    stage2_col18[5] <= stage1_col18[7];
                    stage2_col19[0] <= fa_s1_c18_n17_c;
                    stage2_col19[1] <= fa_s1_c18_n18_c;
                    stage2_col19[2] <= fa_s1_c19_n19_s;
                    stage2_col19[3] <= fa_s1_c19_n20_s;
                    stage2_col19[4] <= stage1_col19[6];
                    stage2_col20[0] <= fa_s1_c19_n19_c;
                    stage2_col20[1] <= fa_s1_c19_n20_c;
                    stage2_col20[2] <= fa_s1_c20_n21_s;
                    stage2_col20[3] <= fa_s1_c20_n22_s;
                    stage2_col20[4] <= stage1_col20[6];
                    stage2_col21[0] <= fa_s1_c20_n21_c;
                    stage2_col21[1] <= fa_s1_c20_n22_c;
                    stage2_col21[2] <= fa_s1_c21_n23_s;
                    stage2_col21[3] <= fa_s1_c21_n24_s;
                    stage2_col21[4] <= fa_s1_c21_n25_s;
                    stage2_col22[0] <= fa_s1_c21_n23_c;
                    stage2_col22[1] <= fa_s1_c21_n24_c;
                    stage2_col22[2] <= fa_s1_c21_n25_c;
                    stage2_col22[3] <= fa_s1_c22_n26_s;
                    stage2_col22[4] <= fa_s1_c22_n27_s;
                    stage2_col22[5] <= stage1_col22[6];
                    stage2_col22[6] <= stage1_col22[7];
                    stage2_col23[0] <= fa_s1_c22_n26_c;
                    stage2_col23[1] <= fa_s1_c22_n27_c;
                    stage2_col23[2] <= fa_s1_c23_n28_s;
                    stage2_col23[3] <= fa_s1_c23_n29_s;
                    stage2_col23[4] <= stage1_col23[6];
                    stage2_col23[5] <= stage1_col23[7];
                    stage2_col24[0] <= fa_s1_c23_n28_c;
                    stage2_col24[1] <= fa_s1_c23_n29_c;
                    stage2_col24[2] <= fa_s1_c24_n30_s;
                    stage2_col24[3] <= fa_s1_c24_n31_s;
                    stage2_col24[4] <= fa_s1_c24_n32_s;
                    stage2_col24[5] <= stage1_col24[9];
                    stage2_col25[0] <= fa_s1_c24_n30_c;
                    stage2_col25[1] <= fa_s1_c24_n31_c;
                    stage2_col25[2] <= fa_s1_c24_n32_c;
                    stage2_col25[3] <= fa_s1_c25_n33_s;
                    stage2_col25[4] <= fa_s1_c25_n34_s;
                    stage2_col25[5] <= fa_s1_c25_n35_s;
                    stage2_col26[0] <= fa_s1_c25_n33_c;
                    stage2_col26[1] <= fa_s1_c25_n34_c;
                    stage2_col26[2] <= fa_s1_c25_n35_c;
                    stage2_col26[3] <= fa_s1_c26_n36_s;
                    stage2_col26[4] <= fa_s1_c26_n37_s;
                    stage2_col26[5] <= fa_s1_c26_n38_s;
                    stage2_col27[0] <= fa_s1_c26_n36_c;
                    stage2_col27[1] <= fa_s1_c26_n37_c;
                    stage2_col27[2] <= fa_s1_c26_n38_c;
                    stage2_col27[3] <= fa_s1_c27_n39_s;
                    stage2_col27[4] <= fa_s1_c27_n40_s;
                    stage2_col27[5] <= fa_s1_c27_n41_s;
                    stage2_col27[6] <= stage1_col27[9];
                    stage2_col27[7] <= stage1_col27[10];
                    stage2_col28[0] <= fa_s1_c27_n39_c;
                    stage2_col28[1] <= fa_s1_c27_n40_c;
                    stage2_col28[2] <= fa_s1_c27_n41_c;
                    stage2_col28[3] <= fa_s1_c28_n42_s;
                    stage2_col28[4] <= fa_s1_c28_n43_s;
                    stage2_col28[5] <= fa_s1_c28_n44_s;
                    stage2_col28[6] <= stage1_col28[9];
                    stage2_col29[0] <= fa_s1_c28_n42_c;
                    stage2_col29[1] <= fa_s1_c28_n43_c;
                    stage2_col29[2] <= fa_s1_c28_n44_c;
                    stage2_col29[3] <= fa_s1_c29_n45_s;
                    stage2_col29[4] <= fa_s1_c29_n46_s;
                    stage2_col29[5] <= fa_s1_c29_n47_s;
                    stage2_col29[6] <= stage1_col29[9];
                    stage2_col30[0] <= fa_s1_c29_n45_c;
                    stage2_col30[1] <= fa_s1_c29_n46_c;
                    stage2_col30[2] <= fa_s1_c29_n47_c;
                    stage2_col30[3] <= fa_s1_c30_n48_s;
                    stage2_col30[4] <= fa_s1_c30_n49_s;
                    stage2_col30[5] <= fa_s1_c30_n50_s;
                    stage2_col30[6] <= fa_s1_c30_n51_s;
                    stage2_col31[0] <= fa_s1_c30_n48_c;
                    stage2_col31[1] <= fa_s1_c30_n49_c;
                    stage2_col31[2] <= fa_s1_c30_n50_c;
                    stage2_col31[3] <= fa_s1_c30_n51_c;
                    stage2_col31[4] <= fa_s1_c31_n52_s;
                    stage2_col31[5] <= fa_s1_c31_n53_s;
                    stage2_col31[6] <= fa_s1_c31_n54_s;
                    stage2_col31[7] <= stage1_col31[9];
                    stage2_col31[8] <= stage1_col31[10];
                    stage2_col32[0] <= fa_s1_c31_n52_c;
                    stage2_col32[1] <= fa_s1_c31_n53_c;
                    stage2_col32[2] <= fa_s1_c31_n54_c;
                    stage2_col32[3] <= fa_s1_c32_n55_s;
                    stage2_col32[4] <= fa_s1_c32_n56_s;
                    stage2_col32[5] <= fa_s1_c32_n57_s;
                    stage2_col32[6] <= stage1_col32[9];
                    stage2_col32[7] <= stage1_col32[10];
                    stage2_col33[0] <= fa_s1_c32_n55_c;
                    stage2_col33[1] <= fa_s1_c32_n56_c;
                    stage2_col33[2] <= fa_s1_c32_n57_c;
                    stage2_col33[3] <= fa_s1_c33_n58_s;
                    stage2_col33[4] <= fa_s1_c33_n59_s;
                    stage2_col33[5] <= fa_s1_c33_n60_s;
                    stage2_col33[6] <= fa_s1_c33_n61_s;
                    stage2_col33[7] <= stage1_col33[12];
                    stage2_col34[0] <= fa_s1_c33_n58_c;
                    stage2_col34[1] <= fa_s1_c33_n59_c;
                    stage2_col34[2] <= fa_s1_c33_n60_c;
                    stage2_col34[3] <= fa_s1_c33_n61_c;
                    stage2_col34[4] <= fa_s1_c34_n62_s;
                    stage2_col34[5] <= fa_s1_c34_n63_s;
                    stage2_col34[6] <= fa_s1_c34_n64_s;
                    stage2_col34[7] <= fa_s1_c34_n65_s;
                    stage2_col35[0] <= fa_s1_c34_n62_c;
                    stage2_col35[1] <= fa_s1_c34_n63_c;
                    stage2_col35[2] <= fa_s1_c34_n64_c;
                    stage2_col35[3] <= fa_s1_c34_n65_c;
                    stage2_col35[4] <= fa_s1_c35_n66_s;
                    stage2_col35[5] <= fa_s1_c35_n67_s;
                    stage2_col35[6] <= fa_s1_c35_n68_s;
                    stage2_col35[7] <= fa_s1_c35_n69_s;
                    stage2_col36[0] <= fa_s1_c35_n66_c;
                    stage2_col36[1] <= fa_s1_c35_n67_c;
                    stage2_col36[2] <= fa_s1_c35_n68_c;
                    stage2_col36[3] <= fa_s1_c35_n69_c;
                    stage2_col36[4] <= fa_s1_c36_n70_s;
                    stage2_col36[5] <= fa_s1_c36_n71_s;
                    stage2_col36[6] <= fa_s1_c36_n72_s;
                    stage2_col36[7] <= fa_s1_c36_n73_s;
                    stage2_col36[8] <= stage1_col36[12];
                    stage2_col36[9] <= stage1_col36[13];
                    stage2_col37[0] <= fa_s1_c36_n70_c;
                    stage2_col37[1] <= fa_s1_c36_n71_c;
                    stage2_col37[2] <= fa_s1_c36_n72_c;
                    stage2_col37[3] <= fa_s1_c36_n73_c;
                    stage2_col37[4] <= fa_s1_c37_n74_s;
                    stage2_col37[5] <= fa_s1_c37_n75_s;
                    stage2_col37[6] <= fa_s1_c37_n76_s;
                    stage2_col37[7] <= fa_s1_c37_n77_s;
                    stage2_col37[8] <= stage1_col37[12];
                    stage2_col38[0] <= fa_s1_c37_n74_c;
                    stage2_col38[1] <= fa_s1_c37_n75_c;
                    stage2_col38[2] <= fa_s1_c37_n76_c;
                    stage2_col38[3] <= fa_s1_c37_n77_c;
                    stage2_col38[4] <= fa_s1_c38_n78_s;
                    stage2_col38[5] <= fa_s1_c38_n79_s;
                    stage2_col38[6] <= fa_s1_c38_n80_s;
                    stage2_col38[7] <= fa_s1_c38_n81_s;
                    stage2_col38[8] <= stage1_col38[12];
                    stage2_col39[0] <= fa_s1_c38_n78_c;
                    stage2_col39[1] <= fa_s1_c38_n79_c;
                    stage2_col39[2] <= fa_s1_c38_n80_c;
                    stage2_col39[3] <= fa_s1_c38_n81_c;
                    stage2_col39[4] <= fa_s1_c39_n82_s;
                    stage2_col39[5] <= fa_s1_c39_n83_s;
                    stage2_col39[6] <= fa_s1_c39_n84_s;
                    stage2_col39[7] <= fa_s1_c39_n85_s;
                    stage2_col39[8] <= fa_s1_c39_n86_s;
                    stage2_col40[0] <= fa_s1_c39_n82_c;
                    stage2_col40[1] <= fa_s1_c39_n83_c;
                    stage2_col40[2] <= fa_s1_c39_n84_c;
                    stage2_col40[3] <= fa_s1_c39_n85_c;
                    stage2_col40[4] <= fa_s1_c39_n86_c;
                    stage2_col40[5] <= fa_s1_c40_n87_s;
                    stage2_col40[6] <= fa_s1_c40_n88_s;
                    stage2_col40[7] <= fa_s1_c40_n89_s;
                    stage2_col40[8] <= fa_s1_c40_n90_s;
                    stage2_col40[9] <= stage1_col40[12];
                    stage2_col40[10] <= stage1_col40[13];
                    stage2_col41[0] <= fa_s1_c40_n87_c;
                    stage2_col41[1] <= fa_s1_c40_n88_c;
                    stage2_col41[2] <= fa_s1_c40_n89_c;
                    stage2_col41[3] <= fa_s1_c40_n90_c;
                    stage2_col41[4] <= fa_s1_c41_n91_s;
                    stage2_col41[5] <= fa_s1_c41_n92_s;
                    stage2_col41[6] <= fa_s1_c41_n93_s;
                    stage2_col41[7] <= fa_s1_c41_n94_s;
                    stage2_col41[8] <= stage1_col41[12];
                    stage2_col41[9] <= stage1_col41[13];
                    stage2_col42[0] <= fa_s1_c41_n91_c;
                    stage2_col42[1] <= fa_s1_c41_n92_c;
                    stage2_col42[2] <= fa_s1_c41_n93_c;
                    stage2_col42[3] <= fa_s1_c41_n94_c;
                    stage2_col42[4] <= fa_s1_c42_n95_s;
                    stage2_col42[5] <= fa_s1_c42_n96_s;
                    stage2_col42[6] <= fa_s1_c42_n97_s;
                    stage2_col42[7] <= fa_s1_c42_n98_s;
                    stage2_col42[8] <= fa_s1_c42_n99_s;
                    stage2_col42[9] <= stage1_col42[15];
                    stage2_col43[0] <= fa_s1_c42_n95_c;
                    stage2_col43[1] <= fa_s1_c42_n96_c;
                    stage2_col43[2] <= fa_s1_c42_n97_c;
                    stage2_col43[3] <= fa_s1_c42_n98_c;
                    stage2_col43[4] <= fa_s1_c42_n99_c;
                    stage2_col43[5] <= fa_s1_c43_n100_s;
                    stage2_col43[6] <= fa_s1_c43_n101_s;
                    stage2_col43[7] <= fa_s1_c43_n102_s;
                    stage2_col43[8] <= fa_s1_c43_n103_s;
                    stage2_col43[9] <= fa_s1_c43_n104_s;
                    stage2_col44[0] <= fa_s1_c43_n100_c;
                    stage2_col44[1] <= fa_s1_c43_n101_c;
                    stage2_col44[2] <= fa_s1_c43_n102_c;
                    stage2_col44[3] <= fa_s1_c43_n103_c;
                    stage2_col44[4] <= fa_s1_c43_n104_c;
                    stage2_col44[5] <= fa_s1_c44_n105_s;
                    stage2_col44[6] <= fa_s1_c44_n106_s;
                    stage2_col44[7] <= fa_s1_c44_n107_s;
                    stage2_col44[8] <= fa_s1_c44_n108_s;
                    stage2_col44[9] <= fa_s1_c44_n109_s;
                    stage2_col45[0] <= fa_s1_c44_n105_c;
                    stage2_col45[1] <= fa_s1_c44_n106_c;
                    stage2_col45[2] <= fa_s1_c44_n107_c;
                    stage2_col45[3] <= fa_s1_c44_n108_c;
                    stage2_col45[4] <= fa_s1_c44_n109_c;
                    stage2_col45[5] <= fa_s1_c45_n110_s;
                    stage2_col45[6] <= fa_s1_c45_n111_s;
                    stage2_col45[7] <= fa_s1_c45_n112_s;
                    stage2_col45[8] <= fa_s1_c45_n113_s;
                    stage2_col45[9] <= fa_s1_c45_n114_s;
                    stage2_col45[10] <= stage1_col45[15];
                    stage2_col45[11] <= stage1_col45[16];
                    stage2_col46[0] <= fa_s1_c45_n110_c;
                    stage2_col46[1] <= fa_s1_c45_n111_c;
                    stage2_col46[2] <= fa_s1_c45_n112_c;
                    stage2_col46[3] <= fa_s1_c45_n113_c;
                    stage2_col46[4] <= fa_s1_c45_n114_c;
                    stage2_col46[5] <= fa_s1_c46_n115_s;
                    stage2_col46[6] <= fa_s1_c46_n116_s;
                    stage2_col46[7] <= fa_s1_c46_n117_s;
                    stage2_col46[8] <= fa_s1_c46_n118_s;
                    stage2_col46[9] <= fa_s1_c46_n119_s;
                    stage2_col46[10] <= stage1_col46[15];
                    stage2_col47[0] <= fa_s1_c46_n115_c;
                    stage2_col47[1] <= fa_s1_c46_n116_c;
                    stage2_col47[2] <= fa_s1_c46_n117_c;
                    stage2_col47[3] <= fa_s1_c46_n118_c;
                    stage2_col47[4] <= fa_s1_c46_n119_c;
                    stage2_col47[5] <= fa_s1_c47_n120_s;
                    stage2_col47[6] <= fa_s1_c47_n121_s;
                    stage2_col47[7] <= fa_s1_c47_n122_s;
                    stage2_col47[8] <= fa_s1_c47_n123_s;
                    stage2_col47[9] <= fa_s1_c47_n124_s;
                    stage2_col47[10] <= stage1_col47[15];
                    stage2_col48[0] <= fa_s1_c47_n120_c;
                    stage2_col48[1] <= fa_s1_c47_n121_c;
                    stage2_col48[2] <= fa_s1_c47_n122_c;
                    stage2_col48[3] <= fa_s1_c47_n123_c;
                    stage2_col48[4] <= fa_s1_c47_n124_c;
                    stage2_col48[5] <= fa_s1_c48_n125_s;
                    stage2_col48[6] <= fa_s1_c48_n126_s;
                    stage2_col48[7] <= fa_s1_c48_n127_s;
                    stage2_col48[8] <= fa_s1_c48_n128_s;
                    stage2_col48[9] <= fa_s1_c48_n129_s;
                    stage2_col48[10] <= fa_s1_c48_n130_s;
                    stage2_col49[0] <= fa_s1_c48_n125_c;
                    stage2_col49[1] <= fa_s1_c48_n126_c;
                    stage2_col49[2] <= fa_s1_c48_n127_c;
                    stage2_col49[3] <= fa_s1_c48_n128_c;
                    stage2_col49[4] <= fa_s1_c48_n129_c;
                    stage2_col49[5] <= fa_s1_c48_n130_c;
                    stage2_col49[6] <= fa_s1_c49_n131_s;
                    stage2_col49[7] <= fa_s1_c49_n132_s;
                    stage2_col49[8] <= fa_s1_c49_n133_s;
                    stage2_col49[9] <= fa_s1_c49_n134_s;
                    stage2_col49[10] <= fa_s1_c49_n135_s;
                    stage2_col49[11] <= stage1_col49[15];
                    stage2_col49[12] <= stage1_col49[16];
                    stage2_col50[0] <= fa_s1_c49_n131_c;
                    stage2_col50[1] <= fa_s1_c49_n132_c;
                    stage2_col50[2] <= fa_s1_c49_n133_c;
                    stage2_col50[3] <= fa_s1_c49_n134_c;
                    stage2_col50[4] <= fa_s1_c49_n135_c;
                    stage2_col50[5] <= fa_s1_c50_n136_s;
                    stage2_col50[6] <= fa_s1_c50_n137_s;
                    stage2_col50[7] <= fa_s1_c50_n138_s;
                    stage2_col50[8] <= fa_s1_c50_n139_s;
                    stage2_col50[9] <= fa_s1_c50_n140_s;
                    stage2_col50[10] <= stage1_col50[15];
                    stage2_col50[11] <= stage1_col50[16];
                    stage2_col51[0] <= fa_s1_c50_n136_c;
                    stage2_col51[1] <= fa_s1_c50_n137_c;
                    stage2_col51[2] <= fa_s1_c50_n138_c;
                    stage2_col51[3] <= fa_s1_c50_n139_c;
                    stage2_col51[4] <= fa_s1_c50_n140_c;
                    stage2_col51[5] <= fa_s1_c51_n141_s;
                    stage2_col51[6] <= fa_s1_c51_n142_s;
                    stage2_col51[7] <= fa_s1_c51_n143_s;
                    stage2_col51[8] <= fa_s1_c51_n144_s;
                    stage2_col51[9] <= fa_s1_c51_n145_s;
                    stage2_col51[10] <= fa_s1_c51_n146_s;
                    stage2_col51[11] <= stage1_col51[18];
                    stage2_col52[0] <= fa_s1_c51_n141_c;
                    stage2_col52[1] <= fa_s1_c51_n142_c;
                    stage2_col52[2] <= fa_s1_c51_n143_c;
                    stage2_col52[3] <= fa_s1_c51_n144_c;
                    stage2_col52[4] <= fa_s1_c51_n145_c;
                    stage2_col52[5] <= fa_s1_c51_n146_c;
                    stage2_col52[6] <= fa_s1_c52_n147_s;
                    stage2_col52[7] <= fa_s1_c52_n148_s;
                    stage2_col52[8] <= fa_s1_c52_n149_s;
                    stage2_col52[9] <= fa_s1_c52_n150_s;
                    stage2_col52[10] <= fa_s1_c52_n151_s;
                    stage2_col52[11] <= fa_s1_c52_n152_s;
                    stage2_col53[0] <= fa_s1_c52_n147_c;
                    stage2_col53[1] <= fa_s1_c52_n148_c;
                    stage2_col53[2] <= fa_s1_c52_n149_c;
                    stage2_col53[3] <= fa_s1_c52_n150_c;
                    stage2_col53[4] <= fa_s1_c52_n151_c;
                    stage2_col53[5] <= fa_s1_c52_n152_c;
                    stage2_col53[6] <= fa_s1_c53_n153_s;
                    stage2_col53[7] <= fa_s1_c53_n154_s;
                    stage2_col53[8] <= fa_s1_c53_n155_s;
                    stage2_col53[9] <= fa_s1_c53_n156_s;
                    stage2_col53[10] <= fa_s1_c53_n157_s;
                    stage2_col53[11] <= fa_s1_c53_n158_s;
                    stage2_col54[0] <= fa_s1_c53_n153_c;
                    stage2_col54[1] <= fa_s1_c53_n154_c;
                    stage2_col54[2] <= fa_s1_c53_n155_c;
                    stage2_col54[3] <= fa_s1_c53_n156_c;
                    stage2_col54[4] <= fa_s1_c53_n157_c;
                    stage2_col54[5] <= fa_s1_c53_n158_c;
                    stage2_col54[6] <= fa_s1_c54_n159_s;
                    stage2_col54[7] <= fa_s1_c54_n160_s;
                    stage2_col54[8] <= fa_s1_c54_n161_s;
                    stage2_col54[9] <= fa_s1_c54_n162_s;
                    stage2_col54[10] <= fa_s1_c54_n163_s;
                    stage2_col54[11] <= fa_s1_c54_n164_s;
                    stage2_col54[12] <= stage1_col54[18];
                    stage2_col54[13] <= stage1_col54[19];
                    stage2_col55[0] <= fa_s1_c54_n159_c;
                    stage2_col55[1] <= fa_s1_c54_n160_c;
                    stage2_col55[2] <= fa_s1_c54_n161_c;
                    stage2_col55[3] <= fa_s1_c54_n162_c;
                    stage2_col55[4] <= fa_s1_c54_n163_c;
                    stage2_col55[5] <= fa_s1_c54_n164_c;
                    stage2_col55[6] <= fa_s1_c55_n165_s;
                    stage2_col55[7] <= fa_s1_c55_n166_s;
                    stage2_col55[8] <= fa_s1_c55_n167_s;
                    stage2_col55[9] <= fa_s1_c55_n168_s;
                    stage2_col55[10] <= fa_s1_c55_n169_s;
                    stage2_col55[11] <= fa_s1_c55_n170_s;
                    stage2_col55[12] <= stage1_col55[18];
                    stage2_col56[0] <= fa_s1_c55_n165_c;
                    stage2_col56[1] <= fa_s1_c55_n166_c;
                    stage2_col56[2] <= fa_s1_c55_n167_c;
                    stage2_col56[3] <= fa_s1_c55_n168_c;
                    stage2_col56[4] <= fa_s1_c55_n169_c;
                    stage2_col56[5] <= fa_s1_c55_n170_c;
                    stage2_col56[6] <= fa_s1_c56_n171_s;
                    stage2_col56[7] <= fa_s1_c56_n172_s;
                    stage2_col56[8] <= fa_s1_c56_n173_s;
                    stage2_col56[9] <= fa_s1_c56_n174_s;
                    stage2_col56[10] <= fa_s1_c56_n175_s;
                    stage2_col56[11] <= fa_s1_c56_n176_s;
                    stage2_col56[12] <= stage1_col56[18];
                    stage2_col57[0] <= fa_s1_c56_n171_c;
                    stage2_col57[1] <= fa_s1_c56_n172_c;
                    stage2_col57[2] <= fa_s1_c56_n173_c;
                    stage2_col57[3] <= fa_s1_c56_n174_c;
                    stage2_col57[4] <= fa_s1_c56_n175_c;
                    stage2_col57[5] <= fa_s1_c56_n176_c;
                    stage2_col57[6] <= fa_s1_c57_n177_s;
                    stage2_col57[7] <= fa_s1_c57_n178_s;
                    stage2_col57[8] <= fa_s1_c57_n179_s;
                    stage2_col57[9] <= fa_s1_c57_n180_s;
                    stage2_col57[10] <= fa_s1_c57_n181_s;
                    stage2_col57[11] <= fa_s1_c57_n182_s;
                    stage2_col57[12] <= fa_s1_c57_n183_s;
                    stage2_col58[0] <= fa_s1_c57_n177_c;
                    stage2_col58[1] <= fa_s1_c57_n178_c;
                    stage2_col58[2] <= fa_s1_c57_n179_c;
                    stage2_col58[3] <= fa_s1_c57_n180_c;
                    stage2_col58[4] <= fa_s1_c57_n181_c;
                    stage2_col58[5] <= fa_s1_c57_n182_c;
                    stage2_col58[6] <= fa_s1_c57_n183_c;
                    stage2_col58[7] <= fa_s1_c58_n184_s;
                    stage2_col58[8] <= fa_s1_c58_n185_s;
                    stage2_col58[9] <= fa_s1_c58_n186_s;
                    stage2_col58[10] <= fa_s1_c58_n187_s;
                    stage2_col58[11] <= fa_s1_c58_n188_s;
                    stage2_col58[12] <= fa_s1_c58_n189_s;
                    stage2_col58[13] <= stage1_col58[18];
                    stage2_col58[14] <= stage1_col58[19];
                    stage2_col59[0] <= fa_s1_c58_n184_c;
                    stage2_col59[1] <= fa_s1_c58_n185_c;
                    stage2_col59[2] <= fa_s1_c58_n186_c;
                    stage2_col59[3] <= fa_s1_c58_n187_c;
                    stage2_col59[4] <= fa_s1_c58_n188_c;
                    stage2_col59[5] <= fa_s1_c58_n189_c;
                    stage2_col59[6] <= fa_s1_c59_n190_s;
                    stage2_col59[7] <= fa_s1_c59_n191_s;
                    stage2_col59[8] <= fa_s1_c59_n192_s;
                    stage2_col59[9] <= fa_s1_c59_n193_s;
                    stage2_col59[10] <= fa_s1_c59_n194_s;
                    stage2_col59[11] <= fa_s1_c59_n195_s;
                    stage2_col59[12] <= stage1_col59[18];
                    stage2_col59[13] <= stage1_col59[19];
                    stage2_col60[0] <= fa_s1_c59_n190_c;
                    stage2_col60[1] <= fa_s1_c59_n191_c;
                    stage2_col60[2] <= fa_s1_c59_n192_c;
                    stage2_col60[3] <= fa_s1_c59_n193_c;
                    stage2_col60[4] <= fa_s1_c59_n194_c;
                    stage2_col60[5] <= fa_s1_c59_n195_c;
                    stage2_col60[6] <= fa_s1_c60_n196_s;
                    stage2_col60[7] <= fa_s1_c60_n197_s;
                    stage2_col60[8] <= fa_s1_c60_n198_s;
                    stage2_col60[9] <= fa_s1_c60_n199_s;
                    stage2_col60[10] <= fa_s1_c60_n200_s;
                    stage2_col60[11] <= fa_s1_c60_n201_s;
                    stage2_col60[12] <= fa_s1_c60_n202_s;
                    stage2_col60[13] <= stage1_col60[21];
                    stage2_col61[0] <= fa_s1_c60_n196_c;
                    stage2_col61[1] <= fa_s1_c60_n197_c;
                    stage2_col61[2] <= fa_s1_c60_n198_c;
                    stage2_col61[3] <= fa_s1_c60_n199_c;
                    stage2_col61[4] <= fa_s1_c60_n200_c;
                    stage2_col61[5] <= fa_s1_c60_n201_c;
                    stage2_col61[6] <= fa_s1_c60_n202_c;
                    stage2_col61[7] <= fa_s1_c61_n203_s;
                    stage2_col61[8] <= fa_s1_c61_n204_s;
                    stage2_col61[9] <= fa_s1_c61_n205_s;
                    stage2_col61[10] <= fa_s1_c61_n206_s;
                    stage2_col61[11] <= fa_s1_c61_n207_s;
                    stage2_col61[12] <= fa_s1_c61_n208_s;
                    stage2_col61[13] <= fa_s1_c61_n209_s;
                    stage2_col62[0] <= fa_s1_c61_n203_c;
                    stage2_col62[1] <= fa_s1_c61_n204_c;
                    stage2_col62[2] <= fa_s1_c61_n205_c;
                    stage2_col62[3] <= fa_s1_c61_n206_c;
                    stage2_col62[4] <= fa_s1_c61_n207_c;
                    stage2_col62[5] <= fa_s1_c61_n208_c;
                    stage2_col62[6] <= fa_s1_c61_n209_c;
                    stage2_col62[7] <= fa_s1_c62_n210_s;
                    stage2_col62[8] <= fa_s1_c62_n211_s;
                    stage2_col62[9] <= fa_s1_c62_n212_s;
                    stage2_col62[10] <= fa_s1_c62_n213_s;
                    stage2_col62[11] <= fa_s1_c62_n214_s;
                    stage2_col62[12] <= fa_s1_c62_n215_s;
                    stage2_col62[13] <= fa_s1_c62_n216_s;
                    stage2_col63[0] <= fa_s1_c62_n210_c;
                    stage2_col63[1] <= fa_s1_c62_n211_c;
                    stage2_col63[2] <= fa_s1_c62_n212_c;
                    stage2_col63[3] <= fa_s1_c62_n213_c;
                    stage2_col63[4] <= fa_s1_c62_n214_c;
                    stage2_col63[5] <= fa_s1_c62_n215_c;
                    stage2_col63[6] <= fa_s1_c62_n216_c;
                    stage2_col63[7] <= fa_s1_c63_n217_s;
                    stage2_col63[8] <= fa_s1_c63_n218_s;
                    stage2_col63[9] <= fa_s1_c63_n219_s;
                    stage2_col63[10] <= fa_s1_c63_n220_s;
                    stage2_col63[11] <= fa_s1_c63_n221_s;
                    stage2_col63[12] <= fa_s1_c63_n222_s;
                    stage2_col63[13] <= fa_s1_c63_n223_s;
                    stage2_col63[14] <= stage1_col63[21];
                    stage2_col63[15] <= stage1_col63[22];
                    stage2_col64[0] <= fa_s1_c63_n217_c;
                    stage2_col64[1] <= fa_s1_c63_n218_c;
                    stage2_col64[2] <= fa_s1_c63_n219_c;
                    stage2_col64[3] <= fa_s1_c63_n220_c;
                    stage2_col64[4] <= fa_s1_c63_n221_c;
                    stage2_col64[5] <= fa_s1_c63_n222_c;
                    stage2_col64[6] <= fa_s1_c63_n223_c;
                    stage2_col64[7] <= fa_s1_c64_n224_s;
                    stage2_col64[8] <= fa_s1_c64_n225_s;
                    stage2_col64[9] <= fa_s1_c64_n226_s;
                    stage2_col64[10] <= fa_s1_c64_n227_s;
                    stage2_col64[11] <= fa_s1_c64_n228_s;
                    stage2_col64[12] <= fa_s1_c64_n229_s;
                    stage2_col64[13] <= fa_s1_c64_n230_s;
                    stage2_col65[0] <= fa_s1_c64_n224_c;
                    stage2_col65[1] <= fa_s1_c64_n225_c;
                    stage2_col65[2] <= fa_s1_c64_n226_c;
                    stage2_col65[3] <= fa_s1_c64_n227_c;
                    stage2_col65[4] <= fa_s1_c64_n228_c;
                    stage2_col65[5] <= fa_s1_c64_n229_c;
                    stage2_col65[6] <= fa_s1_c64_n230_c;
                    stage2_col65[7] <= fa_s1_c65_n231_s;
                    stage2_col65[8] <= fa_s1_c65_n232_s;
                    stage2_col65[9] <= fa_s1_c65_n233_s;
                    stage2_col65[10] <= fa_s1_c65_n234_s;
                    stage2_col65[11] <= fa_s1_c65_n235_s;
                    stage2_col65[12] <= fa_s1_c65_n236_s;
                    stage2_col65[13] <= fa_s1_c65_n237_s;
                    stage2_col65[14] <= stage1_col65[21];
                    stage2_col65[15] <= stage1_col65[22];
                    stage2_col66[0] <= fa_s1_c65_n231_c;
                    stage2_col66[1] <= fa_s1_c65_n232_c;
                    stage2_col66[2] <= fa_s1_c65_n233_c;
                    stage2_col66[3] <= fa_s1_c65_n234_c;
                    stage2_col66[4] <= fa_s1_c65_n235_c;
                    stage2_col66[5] <= fa_s1_c65_n236_c;
                    stage2_col66[6] <= fa_s1_c65_n237_c;
                    stage2_col66[7] <= fa_s1_c66_n238_s;
                    stage2_col66[8] <= fa_s1_c66_n239_s;
                    stage2_col66[9] <= fa_s1_c66_n240_s;
                    stage2_col66[10] <= fa_s1_c66_n241_s;
                    stage2_col66[11] <= fa_s1_c66_n242_s;
                    stage2_col66[12] <= fa_s1_c66_n243_s;
                    stage2_col66[13] <= fa_s1_c66_n244_s;
                    stage2_col67[0] <= fa_s1_c66_n238_c;
                    stage2_col67[1] <= fa_s1_c66_n239_c;
                    stage2_col67[2] <= fa_s1_c66_n240_c;
                    stage2_col67[3] <= fa_s1_c66_n241_c;
                    stage2_col67[4] <= fa_s1_c66_n242_c;
                    stage2_col67[5] <= fa_s1_c66_n243_c;
                    stage2_col67[6] <= fa_s1_c66_n244_c;
                    stage2_col67[7] <= fa_s1_c67_n245_s;
                    stage2_col67[8] <= fa_s1_c67_n246_s;
                    stage2_col67[9] <= fa_s1_c67_n247_s;
                    stage2_col67[10] <= fa_s1_c67_n248_s;
                    stage2_col67[11] <= fa_s1_c67_n249_s;
                    stage2_col67[12] <= fa_s1_c67_n250_s;
                    stage2_col67[13] <= fa_s1_c67_n251_s;
                    stage2_col67[14] <= stage1_col67[21];
                    stage2_col67[15] <= stage1_col67[22];
                    stage2_col68[0] <= fa_s1_c67_n245_c;
                    stage2_col68[1] <= fa_s1_c67_n246_c;
                    stage2_col68[2] <= fa_s1_c67_n247_c;
                    stage2_col68[3] <= fa_s1_c67_n248_c;
                    stage2_col68[4] <= fa_s1_c67_n249_c;
                    stage2_col68[5] <= fa_s1_c67_n250_c;
                    stage2_col68[6] <= fa_s1_c67_n251_c;
                    stage2_col68[7] <= fa_s1_c68_n252_s;
                    stage2_col68[8] <= fa_s1_c68_n253_s;
                    stage2_col68[9] <= fa_s1_c68_n254_s;
                    stage2_col68[10] <= fa_s1_c68_n255_s;
                    stage2_col68[11] <= fa_s1_c68_n256_s;
                    stage2_col68[12] <= fa_s1_c68_n257_s;
                    stage2_col68[13] <= fa_s1_c68_n258_s;
                    stage2_col69[0] <= fa_s1_c68_n252_c;
                    stage2_col69[1] <= fa_s1_c68_n253_c;
                    stage2_col69[2] <= fa_s1_c68_n254_c;
                    stage2_col69[3] <= fa_s1_c68_n255_c;
                    stage2_col69[4] <= fa_s1_c68_n256_c;
                    stage2_col69[5] <= fa_s1_c68_n257_c;
                    stage2_col69[6] <= fa_s1_c68_n258_c;
                    stage2_col69[7] <= fa_s1_c69_n259_s;
                    stage2_col69[8] <= fa_s1_c69_n260_s;
                    stage2_col69[9] <= fa_s1_c69_n261_s;
                    stage2_col69[10] <= fa_s1_c69_n262_s;
                    stage2_col69[11] <= fa_s1_c69_n263_s;
                    stage2_col69[12] <= fa_s1_c69_n264_s;
                    stage2_col69[13] <= fa_s1_c69_n265_s;
                    stage2_col69[14] <= stage1_col69[21];
                    stage2_col69[15] <= stage1_col69[22];
                    stage2_col70[0] <= fa_s1_c69_n259_c;
                    stage2_col70[1] <= fa_s1_c69_n260_c;
                    stage2_col70[2] <= fa_s1_c69_n261_c;
                    stage2_col70[3] <= fa_s1_c69_n262_c;
                    stage2_col70[4] <= fa_s1_c69_n263_c;
                    stage2_col70[5] <= fa_s1_c69_n264_c;
                    stage2_col70[6] <= fa_s1_c69_n265_c;
                    stage2_col70[7] <= fa_s1_c70_n266_s;
                    stage2_col70[8] <= fa_s1_c70_n267_s;
                    stage2_col70[9] <= fa_s1_c70_n268_s;
                    stage2_col70[10] <= fa_s1_c70_n269_s;
                    stage2_col70[11] <= fa_s1_c70_n270_s;
                    stage2_col70[12] <= fa_s1_c70_n271_s;
                    stage2_col70[13] <= fa_s1_c70_n272_s;
                    stage2_col71[0] <= fa_s1_c70_n266_c;
                    stage2_col71[1] <= fa_s1_c70_n267_c;
                    stage2_col71[2] <= fa_s1_c70_n268_c;
                    stage2_col71[3] <= fa_s1_c70_n269_c;
                    stage2_col71[4] <= fa_s1_c70_n270_c;
                    stage2_col71[5] <= fa_s1_c70_n271_c;
                    stage2_col71[6] <= fa_s1_c70_n272_c;
                    stage2_col71[7] <= fa_s1_c71_n273_s;
                    stage2_col71[8] <= fa_s1_c71_n274_s;
                    stage2_col71[9] <= fa_s1_c71_n275_s;
                    stage2_col71[10] <= fa_s1_c71_n276_s;
                    stage2_col71[11] <= fa_s1_c71_n277_s;
                    stage2_col71[12] <= fa_s1_c71_n278_s;
                    stage2_col71[13] <= fa_s1_c71_n279_s;
                    stage2_col71[14] <= stage1_col71[21];
                    stage2_col71[15] <= stage1_col71[22];
                    stage2_col72[0] <= fa_s1_c71_n273_c;
                    stage2_col72[1] <= fa_s1_c71_n274_c;
                    stage2_col72[2] <= fa_s1_c71_n275_c;
                    stage2_col72[3] <= fa_s1_c71_n276_c;
                    stage2_col72[4] <= fa_s1_c71_n277_c;
                    stage2_col72[5] <= fa_s1_c71_n278_c;
                    stage2_col72[6] <= fa_s1_c71_n279_c;
                    stage2_col72[7] <= fa_s1_c72_n280_s;
                    stage2_col72[8] <= fa_s1_c72_n281_s;
                    stage2_col72[9] <= fa_s1_c72_n282_s;
                    stage2_col72[10] <= fa_s1_c72_n283_s;
                    stage2_col72[11] <= fa_s1_c72_n284_s;
                    stage2_col72[12] <= fa_s1_c72_n285_s;
                    stage2_col72[13] <= fa_s1_c72_n286_s;
                    stage2_col73[0] <= fa_s1_c72_n280_c;
                    stage2_col73[1] <= fa_s1_c72_n281_c;
                    stage2_col73[2] <= fa_s1_c72_n282_c;
                    stage2_col73[3] <= fa_s1_c72_n283_c;
                    stage2_col73[4] <= fa_s1_c72_n284_c;
                    stage2_col73[5] <= fa_s1_c72_n285_c;
                    stage2_col73[6] <= fa_s1_c72_n286_c;
                    stage2_col73[7] <= fa_s1_c73_n287_s;
                    stage2_col73[8] <= fa_s1_c73_n288_s;
                    stage2_col73[9] <= fa_s1_c73_n289_s;
                    stage2_col73[10] <= fa_s1_c73_n290_s;
                    stage2_col73[11] <= fa_s1_c73_n291_s;
                    stage2_col73[12] <= fa_s1_c73_n292_s;
                    stage2_col73[13] <= fa_s1_c73_n293_s;
                    stage2_col73[14] <= stage1_col73[21];
                    stage2_col73[15] <= stage1_col73[22];
                    stage2_col74[0] <= fa_s1_c73_n287_c;
                    stage2_col74[1] <= fa_s1_c73_n288_c;
                    stage2_col74[2] <= fa_s1_c73_n289_c;
                    stage2_col74[3] <= fa_s1_c73_n290_c;
                    stage2_col74[4] <= fa_s1_c73_n291_c;
                    stage2_col74[5] <= fa_s1_c73_n292_c;
                    stage2_col74[6] <= fa_s1_c73_n293_c;
                    stage2_col74[7] <= fa_s1_c74_n294_s;
                    stage2_col74[8] <= fa_s1_c74_n295_s;
                    stage2_col74[9] <= fa_s1_c74_n296_s;
                    stage2_col74[10] <= fa_s1_c74_n297_s;
                    stage2_col74[11] <= fa_s1_c74_n298_s;
                    stage2_col74[12] <= fa_s1_c74_n299_s;
                    stage2_col74[13] <= fa_s1_c74_n300_s;
                    stage2_col75[0] <= fa_s1_c74_n294_c;
                    stage2_col75[1] <= fa_s1_c74_n295_c;
                    stage2_col75[2] <= fa_s1_c74_n296_c;
                    stage2_col75[3] <= fa_s1_c74_n297_c;
                    stage2_col75[4] <= fa_s1_c74_n298_c;
                    stage2_col75[5] <= fa_s1_c74_n299_c;
                    stage2_col75[6] <= fa_s1_c74_n300_c;
                    stage2_col75[7] <= fa_s1_c75_n301_s;
                    stage2_col75[8] <= fa_s1_c75_n302_s;
                    stage2_col75[9] <= fa_s1_c75_n303_s;
                    stage2_col75[10] <= fa_s1_c75_n304_s;
                    stage2_col75[11] <= fa_s1_c75_n305_s;
                    stage2_col75[12] <= fa_s1_c75_n306_s;
                    stage2_col75[13] <= fa_s1_c75_n307_s;
                    stage2_col75[14] <= stage1_col75[21];
                    stage2_col75[15] <= stage1_col75[22];
                    stage2_col76[0] <= fa_s1_c75_n301_c;
                    stage2_col76[1] <= fa_s1_c75_n302_c;
                    stage2_col76[2] <= fa_s1_c75_n303_c;
                    stage2_col76[3] <= fa_s1_c75_n304_c;
                    stage2_col76[4] <= fa_s1_c75_n305_c;
                    stage2_col76[5] <= fa_s1_c75_n306_c;
                    stage2_col76[6] <= fa_s1_c75_n307_c;
                    stage2_col76[7] <= fa_s1_c76_n308_s;
                    stage2_col76[8] <= fa_s1_c76_n309_s;
                    stage2_col76[9] <= fa_s1_c76_n310_s;
                    stage2_col76[10] <= fa_s1_c76_n311_s;
                    stage2_col76[11] <= fa_s1_c76_n312_s;
                    stage2_col76[12] <= fa_s1_c76_n313_s;
                    stage2_col76[13] <= fa_s1_c76_n314_s;
                    stage2_col77[0] <= fa_s1_c76_n308_c;
                    stage2_col77[1] <= fa_s1_c76_n309_c;
                    stage2_col77[2] <= fa_s1_c76_n310_c;
                    stage2_col77[3] <= fa_s1_c76_n311_c;
                    stage2_col77[4] <= fa_s1_c76_n312_c;
                    stage2_col77[5] <= fa_s1_c76_n313_c;
                    stage2_col77[6] <= fa_s1_c76_n314_c;
                    stage2_col77[7] <= fa_s1_c77_n315_s;
                    stage2_col77[8] <= fa_s1_c77_n316_s;
                    stage2_col77[9] <= fa_s1_c77_n317_s;
                    stage2_col77[10] <= fa_s1_c77_n318_s;
                    stage2_col77[11] <= fa_s1_c77_n319_s;
                    stage2_col77[12] <= fa_s1_c77_n320_s;
                    stage2_col77[13] <= fa_s1_c77_n321_s;
                    stage2_col77[14] <= stage1_col77[21];
                    stage2_col77[15] <= stage1_col77[22];
                    stage2_col78[0] <= fa_s1_c77_n315_c;
                    stage2_col78[1] <= fa_s1_c77_n316_c;
                    stage2_col78[2] <= fa_s1_c77_n317_c;
                    stage2_col78[3] <= fa_s1_c77_n318_c;
                    stage2_col78[4] <= fa_s1_c77_n319_c;
                    stage2_col78[5] <= fa_s1_c77_n320_c;
                    stage2_col78[6] <= fa_s1_c77_n321_c;
                    stage2_col78[7] <= fa_s1_c78_n322_s;
                    stage2_col78[8] <= fa_s1_c78_n323_s;
                    stage2_col78[9] <= fa_s1_c78_n324_s;
                    stage2_col78[10] <= fa_s1_c78_n325_s;
                    stage2_col78[11] <= fa_s1_c78_n326_s;
                    stage2_col78[12] <= fa_s1_c78_n327_s;
                    stage2_col78[13] <= fa_s1_c78_n328_s;
                    stage2_col79[0] <= fa_s1_c78_n322_c;
                    stage2_col79[1] <= fa_s1_c78_n323_c;
                    stage2_col79[2] <= fa_s1_c78_n324_c;
                    stage2_col79[3] <= fa_s1_c78_n325_c;
                    stage2_col79[4] <= fa_s1_c78_n326_c;
                    stage2_col79[5] <= fa_s1_c78_n327_c;
                    stage2_col79[6] <= fa_s1_c78_n328_c;
                    stage2_col79[7] <= fa_s1_c79_n329_s;
                    stage2_col79[8] <= fa_s1_c79_n330_s;
                    stage2_col79[9] <= fa_s1_c79_n331_s;
                    stage2_col79[10] <= fa_s1_c79_n332_s;
                    stage2_col79[11] <= fa_s1_c79_n333_s;
                    stage2_col79[12] <= fa_s1_c79_n334_s;
                    stage2_col79[13] <= fa_s1_c79_n335_s;
                    stage2_col79[14] <= stage1_col79[21];
                    stage2_col79[15] <= stage1_col79[22];
                    stage2_col80[0] <= fa_s1_c79_n329_c;
                    stage2_col80[1] <= fa_s1_c79_n330_c;
                    stage2_col80[2] <= fa_s1_c79_n331_c;
                    stage2_col80[3] <= fa_s1_c79_n332_c;
                    stage2_col80[4] <= fa_s1_c79_n333_c;
                    stage2_col80[5] <= fa_s1_c79_n334_c;
                    stage2_col80[6] <= fa_s1_c79_n335_c;
                    stage2_col80[7] <= fa_s1_c80_n336_s;
                    stage2_col80[8] <= fa_s1_c80_n337_s;
                    stage2_col80[9] <= fa_s1_c80_n338_s;
                    stage2_col80[10] <= fa_s1_c80_n339_s;
                    stage2_col80[11] <= fa_s1_c80_n340_s;
                    stage2_col80[12] <= fa_s1_c80_n341_s;
                    stage2_col80[13] <= fa_s1_c80_n342_s;
                    stage2_col81[0] <= fa_s1_c80_n336_c;
                    stage2_col81[1] <= fa_s1_c80_n337_c;
                    stage2_col81[2] <= fa_s1_c80_n338_c;
                    stage2_col81[3] <= fa_s1_c80_n339_c;
                    stage2_col81[4] <= fa_s1_c80_n340_c;
                    stage2_col81[5] <= fa_s1_c80_n341_c;
                    stage2_col81[6] <= fa_s1_c80_n342_c;
                    stage2_col81[7] <= fa_s1_c81_n343_s;
                    stage2_col81[8] <= fa_s1_c81_n344_s;
                    stage2_col81[9] <= fa_s1_c81_n345_s;
                    stage2_col81[10] <= fa_s1_c81_n346_s;
                    stage2_col81[11] <= fa_s1_c81_n347_s;
                    stage2_col81[12] <= fa_s1_c81_n348_s;
                    stage2_col81[13] <= fa_s1_c81_n349_s;
                    stage2_col81[14] <= stage1_col81[21];
                    stage2_col81[15] <= stage1_col81[22];
                    stage2_col82[0] <= fa_s1_c81_n343_c;
                    stage2_col82[1] <= fa_s1_c81_n344_c;
                    stage2_col82[2] <= fa_s1_c81_n345_c;
                    stage2_col82[3] <= fa_s1_c81_n346_c;
                    stage2_col82[4] <= fa_s1_c81_n347_c;
                    stage2_col82[5] <= fa_s1_c81_n348_c;
                    stage2_col82[6] <= fa_s1_c81_n349_c;
                    stage2_col82[7] <= fa_s1_c82_n350_s;
                    stage2_col82[8] <= fa_s1_c82_n351_s;
                    stage2_col82[9] <= fa_s1_c82_n352_s;
                    stage2_col82[10] <= fa_s1_c82_n353_s;
                    stage2_col82[11] <= fa_s1_c82_n354_s;
                    stage2_col82[12] <= fa_s1_c82_n355_s;
                    stage2_col82[13] <= fa_s1_c82_n356_s;
                    stage2_col83[0] <= fa_s1_c82_n350_c;
                    stage2_col83[1] <= fa_s1_c82_n351_c;
                    stage2_col83[2] <= fa_s1_c82_n352_c;
                    stage2_col83[3] <= fa_s1_c82_n353_c;
                    stage2_col83[4] <= fa_s1_c82_n354_c;
                    stage2_col83[5] <= fa_s1_c82_n355_c;
                    stage2_col83[6] <= fa_s1_c82_n356_c;
                    stage2_col83[7] <= fa_s1_c83_n357_s;
                    stage2_col83[8] <= fa_s1_c83_n358_s;
                    stage2_col83[9] <= fa_s1_c83_n359_s;
                    stage2_col83[10] <= fa_s1_c83_n360_s;
                    stage2_col83[11] <= fa_s1_c83_n361_s;
                    stage2_col83[12] <= fa_s1_c83_n362_s;
                    stage2_col83[13] <= fa_s1_c83_n363_s;
                    stage2_col83[14] <= stage1_col83[21];
                    stage2_col83[15] <= stage1_col83[22];
                    stage2_col84[0] <= fa_s1_c83_n357_c;
                    stage2_col84[1] <= fa_s1_c83_n358_c;
                    stage2_col84[2] <= fa_s1_c83_n359_c;
                    stage2_col84[3] <= fa_s1_c83_n360_c;
                    stage2_col84[4] <= fa_s1_c83_n361_c;
                    stage2_col84[5] <= fa_s1_c83_n362_c;
                    stage2_col84[6] <= fa_s1_c83_n363_c;
                    stage2_col84[7] <= fa_s1_c84_n364_s;
                    stage2_col84[8] <= fa_s1_c84_n365_s;
                    stage2_col84[9] <= fa_s1_c84_n366_s;
                    stage2_col84[10] <= fa_s1_c84_n367_s;
                    stage2_col84[11] <= fa_s1_c84_n368_s;
                    stage2_col84[12] <= fa_s1_c84_n369_s;
                    stage2_col84[13] <= fa_s1_c84_n370_s;
                    stage2_col85[0] <= fa_s1_c84_n364_c;
                    stage2_col85[1] <= fa_s1_c84_n365_c;
                    stage2_col85[2] <= fa_s1_c84_n366_c;
                    stage2_col85[3] <= fa_s1_c84_n367_c;
                    stage2_col85[4] <= fa_s1_c84_n368_c;
                    stage2_col85[5] <= fa_s1_c84_n369_c;
                    stage2_col85[6] <= fa_s1_c84_n370_c;
                    stage2_col85[7] <= fa_s1_c85_n371_s;
                    stage2_col85[8] <= fa_s1_c85_n372_s;
                    stage2_col85[9] <= fa_s1_c85_n373_s;
                    stage2_col85[10] <= fa_s1_c85_n374_s;
                    stage2_col85[11] <= fa_s1_c85_n375_s;
                    stage2_col85[12] <= fa_s1_c85_n376_s;
                    stage2_col85[13] <= fa_s1_c85_n377_s;
                    stage2_col85[14] <= stage1_col85[21];
                    stage2_col85[15] <= stage1_col85[22];
                    stage2_col86[0] <= fa_s1_c85_n371_c;
                    stage2_col86[1] <= fa_s1_c85_n372_c;
                    stage2_col86[2] <= fa_s1_c85_n373_c;
                    stage2_col86[3] <= fa_s1_c85_n374_c;
                    stage2_col86[4] <= fa_s1_c85_n375_c;
                    stage2_col86[5] <= fa_s1_c85_n376_c;
                    stage2_col86[6] <= fa_s1_c85_n377_c;
                    stage2_col86[7] <= fa_s1_c86_n378_s;
                    stage2_col86[8] <= fa_s1_c86_n379_s;
                    stage2_col86[9] <= fa_s1_c86_n380_s;
                    stage2_col86[10] <= fa_s1_c86_n381_s;
                    stage2_col86[11] <= fa_s1_c86_n382_s;
                    stage2_col86[12] <= fa_s1_c86_n383_s;
                    stage2_col86[13] <= fa_s1_c86_n384_s;
                    stage2_col87[0] <= fa_s1_c86_n378_c;
                    stage2_col87[1] <= fa_s1_c86_n379_c;
                    stage2_col87[2] <= fa_s1_c86_n380_c;
                    stage2_col87[3] <= fa_s1_c86_n381_c;
                    stage2_col87[4] <= fa_s1_c86_n382_c;
                    stage2_col87[5] <= fa_s1_c86_n383_c;
                    stage2_col87[6] <= fa_s1_c86_n384_c;
                    stage2_col87[7] <= fa_s1_c87_n385_s;
                    stage2_col87[8] <= fa_s1_c87_n386_s;
                    stage2_col87[9] <= fa_s1_c87_n387_s;
                    stage2_col87[10] <= fa_s1_c87_n388_s;
                    stage2_col87[11] <= fa_s1_c87_n389_s;
                    stage2_col87[12] <= fa_s1_c87_n390_s;
                    stage2_col87[13] <= fa_s1_c87_n391_s;
                    stage2_col87[14] <= stage1_col87[21];
                    stage2_col87[15] <= stage1_col87[22];
                    stage2_col88[0] <= fa_s1_c87_n385_c;
                    stage2_col88[1] <= fa_s1_c87_n386_c;
                    stage2_col88[2] <= fa_s1_c87_n387_c;
                    stage2_col88[3] <= fa_s1_c87_n388_c;
                    stage2_col88[4] <= fa_s1_c87_n389_c;
                    stage2_col88[5] <= fa_s1_c87_n390_c;
                    stage2_col88[6] <= fa_s1_c87_n391_c;
                    stage2_col88[7] <= fa_s1_c88_n392_s;
                    stage2_col88[8] <= fa_s1_c88_n393_s;
                    stage2_col88[9] <= fa_s1_c88_n394_s;
                    stage2_col88[10] <= fa_s1_c88_n395_s;
                    stage2_col88[11] <= fa_s1_c88_n396_s;
                    stage2_col88[12] <= fa_s1_c88_n397_s;
                    stage2_col88[13] <= fa_s1_c88_n398_s;
                    stage2_col89[0] <= fa_s1_c88_n392_c;
                    stage2_col89[1] <= fa_s1_c88_n393_c;
                    stage2_col89[2] <= fa_s1_c88_n394_c;
                    stage2_col89[3] <= fa_s1_c88_n395_c;
                    stage2_col89[4] <= fa_s1_c88_n396_c;
                    stage2_col89[5] <= fa_s1_c88_n397_c;
                    stage2_col89[6] <= fa_s1_c88_n398_c;
                    stage2_col89[7] <= fa_s1_c89_n399_s;
                    stage2_col89[8] <= fa_s1_c89_n400_s;
                    stage2_col89[9] <= fa_s1_c89_n401_s;
                    stage2_col89[10] <= fa_s1_c89_n402_s;
                    stage2_col89[11] <= fa_s1_c89_n403_s;
                    stage2_col89[12] <= fa_s1_c89_n404_s;
                    stage2_col89[13] <= fa_s1_c89_n405_s;
                    stage2_col89[14] <= stage1_col89[21];
                    stage2_col89[15] <= stage1_col89[22];
                    stage2_col90[0] <= fa_s1_c89_n399_c;
                    stage2_col90[1] <= fa_s1_c89_n400_c;
                    stage2_col90[2] <= fa_s1_c89_n401_c;
                    stage2_col90[3] <= fa_s1_c89_n402_c;
                    stage2_col90[4] <= fa_s1_c89_n403_c;
                    stage2_col90[5] <= fa_s1_c89_n404_c;
                    stage2_col90[6] <= fa_s1_c89_n405_c;
                    stage2_col90[7] <= fa_s1_c90_n406_s;
                    stage2_col90[8] <= fa_s1_c90_n407_s;
                    stage2_col90[9] <= fa_s1_c90_n408_s;
                    stage2_col90[10] <= fa_s1_c90_n409_s;
                    stage2_col90[11] <= fa_s1_c90_n410_s;
                    stage2_col90[12] <= fa_s1_c90_n411_s;
                    stage2_col90[13] <= fa_s1_c90_n412_s;
                    stage2_col91[0] <= fa_s1_c90_n406_c;
                    stage2_col91[1] <= fa_s1_c90_n407_c;
                    stage2_col91[2] <= fa_s1_c90_n408_c;
                    stage2_col91[3] <= fa_s1_c90_n409_c;
                    stage2_col91[4] <= fa_s1_c90_n410_c;
                    stage2_col91[5] <= fa_s1_c90_n411_c;
                    stage2_col91[6] <= fa_s1_c90_n412_c;
                    stage2_col91[7] <= fa_s1_c91_n413_s;
                    stage2_col91[8] <= fa_s1_c91_n414_s;
                    stage2_col91[9] <= fa_s1_c91_n415_s;
                    stage2_col91[10] <= fa_s1_c91_n416_s;
                    stage2_col91[11] <= fa_s1_c91_n417_s;
                    stage2_col91[12] <= fa_s1_c91_n418_s;
                    stage2_col91[13] <= fa_s1_c91_n419_s;
                    stage2_col91[14] <= stage1_col91[21];
                    stage2_col91[15] <= stage1_col91[22];
                    stage2_col92[0] <= fa_s1_c91_n413_c;
                    stage2_col92[1] <= fa_s1_c91_n414_c;
                    stage2_col92[2] <= fa_s1_c91_n415_c;
                    stage2_col92[3] <= fa_s1_c91_n416_c;
                    stage2_col92[4] <= fa_s1_c91_n417_c;
                    stage2_col92[5] <= fa_s1_c91_n418_c;
                    stage2_col92[6] <= fa_s1_c91_n419_c;
                    stage2_col92[7] <= fa_s1_c92_n420_s;
                    stage2_col92[8] <= fa_s1_c92_n421_s;
                    stage2_col92[9] <= fa_s1_c92_n422_s;
                    stage2_col92[10] <= fa_s1_c92_n423_s;
                    stage2_col92[11] <= fa_s1_c92_n424_s;
                    stage2_col92[12] <= fa_s1_c92_n425_s;
                    stage2_col92[13] <= fa_s1_c92_n426_s;
                    stage2_col93[0] <= fa_s1_c92_n420_c;
                    stage2_col93[1] <= fa_s1_c92_n421_c;
                    stage2_col93[2] <= fa_s1_c92_n422_c;
                    stage2_col93[3] <= fa_s1_c92_n423_c;
                    stage2_col93[4] <= fa_s1_c92_n424_c;
                    stage2_col93[5] <= fa_s1_c92_n425_c;
                    stage2_col93[6] <= fa_s1_c92_n426_c;
                    stage2_col93[7] <= fa_s1_c93_n427_s;
                    stage2_col93[8] <= fa_s1_c93_n428_s;
                    stage2_col93[9] <= fa_s1_c93_n429_s;
                    stage2_col93[10] <= fa_s1_c93_n430_s;
                    stage2_col93[11] <= fa_s1_c93_n431_s;
                    stage2_col93[12] <= fa_s1_c93_n432_s;
                    stage2_col93[13] <= fa_s1_c93_n433_s;
                    stage2_col93[14] <= stage1_col93[21];
                    stage2_col93[15] <= stage1_col93[22];
                    stage2_col94[0] <= fa_s1_c93_n427_c;
                    stage2_col94[1] <= fa_s1_c93_n428_c;
                    stage2_col94[2] <= fa_s1_c93_n429_c;
                    stage2_col94[3] <= fa_s1_c93_n430_c;
                    stage2_col94[4] <= fa_s1_c93_n431_c;
                    stage2_col94[5] <= fa_s1_c93_n432_c;
                    stage2_col94[6] <= fa_s1_c93_n433_c;
                    stage2_col94[7] <= fa_s1_c94_n434_s;
                    stage2_col94[8] <= fa_s1_c94_n435_s;
                    stage2_col94[9] <= fa_s1_c94_n436_s;
                    stage2_col94[10] <= fa_s1_c94_n437_s;
                    stage2_col94[11] <= fa_s1_c94_n438_s;
                    stage2_col94[12] <= fa_s1_c94_n439_s;
                    stage2_col94[13] <= fa_s1_c94_n440_s;
                    stage2_col95[0] <= fa_s1_c94_n434_c;
                    stage2_col95[1] <= fa_s1_c94_n435_c;
                    stage2_col95[2] <= fa_s1_c94_n436_c;
                    stage2_col95[3] <= fa_s1_c94_n437_c;
                    stage2_col95[4] <= fa_s1_c94_n438_c;
                    stage2_col95[5] <= fa_s1_c94_n439_c;
                    stage2_col95[6] <= fa_s1_c94_n440_c;
                    stage2_col95[7] <= fa_s1_c95_n441_s;
                    stage2_col95[8] <= fa_s1_c95_n442_s;
                    stage2_col95[9] <= fa_s1_c95_n443_s;
                    stage2_col95[10] <= fa_s1_c95_n444_s;
                    stage2_col95[11] <= fa_s1_c95_n445_s;
                    stage2_col95[12] <= fa_s1_c95_n446_s;
                    stage2_col95[13] <= fa_s1_c95_n447_s;
                    stage2_col95[14] <= stage1_col95[21];
                    stage2_col95[15] <= stage1_col95[22];
                    stage2_col96[0] <= fa_s1_c95_n441_c;
                    stage2_col96[1] <= fa_s1_c95_n442_c;
                    stage2_col96[2] <= fa_s1_c95_n443_c;
                    stage2_col96[3] <= fa_s1_c95_n444_c;
                    stage2_col96[4] <= fa_s1_c95_n445_c;
                    stage2_col96[5] <= fa_s1_c95_n446_c;
                    stage2_col96[6] <= fa_s1_c95_n447_c;
                    stage2_col96[7] <= fa_s1_c96_n448_s;
                    stage2_col96[8] <= fa_s1_c96_n449_s;
                    stage2_col96[9] <= fa_s1_c96_n450_s;
                    stage2_col96[10] <= fa_s1_c96_n451_s;
                    stage2_col96[11] <= fa_s1_c96_n452_s;
                    stage2_col96[12] <= fa_s1_c96_n453_s;
                    stage2_col96[13] <= fa_s1_c96_n454_s;
                    stage2_col97[0] <= fa_s1_c96_n448_c;
                    stage2_col97[1] <= fa_s1_c96_n449_c;
                    stage2_col97[2] <= fa_s1_c96_n450_c;
                    stage2_col97[3] <= fa_s1_c96_n451_c;
                    stage2_col97[4] <= fa_s1_c96_n452_c;
                    stage2_col97[5] <= fa_s1_c96_n453_c;
                    stage2_col97[6] <= fa_s1_c96_n454_c;
                    stage2_col97[7] <= fa_s1_c97_n455_s;
                    stage2_col97[8] <= fa_s1_c97_n456_s;
                    stage2_col97[9] <= fa_s1_c97_n457_s;
                    stage2_col97[10] <= fa_s1_c97_n458_s;
                    stage2_col97[11] <= fa_s1_c97_n459_s;
                    stage2_col97[12] <= fa_s1_c97_n460_s;
                    stage2_col97[13] <= fa_s1_c97_n461_s;
                    stage2_col97[14] <= stage1_col97[21];
                    stage2_col97[15] <= stage1_col97[22];
                    stage2_col98[0] <= fa_s1_c97_n455_c;
                    stage2_col98[1] <= fa_s1_c97_n456_c;
                    stage2_col98[2] <= fa_s1_c97_n457_c;
                    stage2_col98[3] <= fa_s1_c97_n458_c;
                    stage2_col98[4] <= fa_s1_c97_n459_c;
                    stage2_col98[5] <= fa_s1_c97_n460_c;
                    stage2_col98[6] <= fa_s1_c97_n461_c;
                    stage2_col98[7] <= fa_s1_c98_n462_s;
                    stage2_col98[8] <= fa_s1_c98_n463_s;
                    stage2_col98[9] <= fa_s1_c98_n464_s;
                    stage2_col98[10] <= fa_s1_c98_n465_s;
                    stage2_col98[11] <= fa_s1_c98_n466_s;
                    stage2_col98[12] <= fa_s1_c98_n467_s;
                    stage2_col98[13] <= fa_s1_c98_n468_s;
                    stage2_col99[0] <= fa_s1_c98_n462_c;
                    stage2_col99[1] <= fa_s1_c98_n463_c;
                    stage2_col99[2] <= fa_s1_c98_n464_c;
                    stage2_col99[3] <= fa_s1_c98_n465_c;
                    stage2_col99[4] <= fa_s1_c98_n466_c;
                    stage2_col99[5] <= fa_s1_c98_n467_c;
                    stage2_col99[6] <= fa_s1_c98_n468_c;
                    stage2_col99[7] <= fa_s1_c99_n469_s;
                    stage2_col99[8] <= fa_s1_c99_n470_s;
                    stage2_col99[9] <= fa_s1_c99_n471_s;
                    stage2_col99[10] <= fa_s1_c99_n472_s;
                    stage2_col99[11] <= fa_s1_c99_n473_s;
                    stage2_col99[12] <= fa_s1_c99_n474_s;
                    stage2_col99[13] <= fa_s1_c99_n475_s;
                    stage2_col99[14] <= stage1_col99[21];
                    stage2_col99[15] <= stage1_col99[22];
                    stage2_col100[0] <= fa_s1_c99_n469_c;
                    stage2_col100[1] <= fa_s1_c99_n470_c;
                    stage2_col100[2] <= fa_s1_c99_n471_c;
                    stage2_col100[3] <= fa_s1_c99_n472_c;
                    stage2_col100[4] <= fa_s1_c99_n473_c;
                    stage2_col100[5] <= fa_s1_c99_n474_c;
                    stage2_col100[6] <= fa_s1_c99_n475_c;
                    stage2_col100[7] <= fa_s1_c100_n476_s;
                    stage2_col100[8] <= fa_s1_c100_n477_s;
                    stage2_col100[9] <= fa_s1_c100_n478_s;
                    stage2_col100[10] <= fa_s1_c100_n479_s;
                    stage2_col100[11] <= fa_s1_c100_n480_s;
                    stage2_col100[12] <= fa_s1_c100_n481_s;
                    stage2_col100[13] <= fa_s1_c100_n482_s;
                    stage2_col101[0] <= fa_s1_c100_n476_c;
                    stage2_col101[1] <= fa_s1_c100_n477_c;
                    stage2_col101[2] <= fa_s1_c100_n478_c;
                    stage2_col101[3] <= fa_s1_c100_n479_c;
                    stage2_col101[4] <= fa_s1_c100_n480_c;
                    stage2_col101[5] <= fa_s1_c100_n481_c;
                    stage2_col101[6] <= fa_s1_c100_n482_c;
                    stage2_col101[7] <= fa_s1_c101_n483_s;
                    stage2_col101[8] <= fa_s1_c101_n484_s;
                    stage2_col101[9] <= fa_s1_c101_n485_s;
                    stage2_col101[10] <= fa_s1_c101_n486_s;
                    stage2_col101[11] <= fa_s1_c101_n487_s;
                    stage2_col101[12] <= fa_s1_c101_n488_s;
                    stage2_col101[13] <= fa_s1_c101_n489_s;
                    stage2_col101[14] <= stage1_col101[21];
                    stage2_col101[15] <= stage1_col101[22];
                    stage2_col102[0] <= fa_s1_c101_n483_c;
                    stage2_col102[1] <= fa_s1_c101_n484_c;
                    stage2_col102[2] <= fa_s1_c101_n485_c;
                    stage2_col102[3] <= fa_s1_c101_n486_c;
                    stage2_col102[4] <= fa_s1_c101_n487_c;
                    stage2_col102[5] <= fa_s1_c101_n488_c;
                    stage2_col102[6] <= fa_s1_c101_n489_c;
                    stage2_col102[7] <= fa_s1_c102_n490_s;
                    stage2_col102[8] <= fa_s1_c102_n491_s;
                    stage2_col102[9] <= fa_s1_c102_n492_s;
                    stage2_col102[10] <= fa_s1_c102_n493_s;
                    stage2_col102[11] <= fa_s1_c102_n494_s;
                    stage2_col102[12] <= fa_s1_c102_n495_s;
                    stage2_col102[13] <= fa_s1_c102_n496_s;
                    stage2_col103[0] <= fa_s1_c102_n490_c;
                    stage2_col103[1] <= fa_s1_c102_n491_c;
                    stage2_col103[2] <= fa_s1_c102_n492_c;
                    stage2_col103[3] <= fa_s1_c102_n493_c;
                    stage2_col103[4] <= fa_s1_c102_n494_c;
                    stage2_col103[5] <= fa_s1_c102_n495_c;
                    stage2_col103[6] <= fa_s1_c102_n496_c;
                    stage2_col103[7] <= fa_s1_c103_n497_s;
                    stage2_col103[8] <= fa_s1_c103_n498_s;
                    stage2_col103[9] <= fa_s1_c103_n499_s;
                    stage2_col103[10] <= fa_s1_c103_n500_s;
                    stage2_col103[11] <= fa_s1_c103_n501_s;
                    stage2_col103[12] <= fa_s1_c103_n502_s;
                    stage2_col103[13] <= fa_s1_c103_n503_s;
                    stage2_col103[14] <= stage1_col103[21];
                    stage2_col103[15] <= stage1_col103[22];
                    stage2_col104[0] <= fa_s1_c103_n497_c;
                    stage2_col104[1] <= fa_s1_c103_n498_c;
                    stage2_col104[2] <= fa_s1_c103_n499_c;
                    stage2_col104[3] <= fa_s1_c103_n500_c;
                    stage2_col104[4] <= fa_s1_c103_n501_c;
                    stage2_col104[5] <= fa_s1_c103_n502_c;
                    stage2_col104[6] <= fa_s1_c103_n503_c;
                    stage2_col104[7] <= fa_s1_c104_n504_s;
                    stage2_col104[8] <= fa_s1_c104_n505_s;
                    stage2_col104[9] <= fa_s1_c104_n506_s;
                    stage2_col104[10] <= fa_s1_c104_n507_s;
                    stage2_col104[11] <= fa_s1_c104_n508_s;
                    stage2_col104[12] <= fa_s1_c104_n509_s;
                    stage2_col104[13] <= fa_s1_c104_n510_s;
                    stage2_col105[0] <= fa_s1_c104_n504_c;
                    stage2_col105[1] <= fa_s1_c104_n505_c;
                    stage2_col105[2] <= fa_s1_c104_n506_c;
                    stage2_col105[3] <= fa_s1_c104_n507_c;
                    stage2_col105[4] <= fa_s1_c104_n508_c;
                    stage2_col105[5] <= fa_s1_c104_n509_c;
                    stage2_col105[6] <= fa_s1_c104_n510_c;
                    stage2_col105[7] <= fa_s1_c105_n511_s;
                    stage2_col105[8] <= fa_s1_c105_n512_s;
                    stage2_col105[9] <= fa_s1_c105_n513_s;
                    stage2_col105[10] <= fa_s1_c105_n514_s;
                    stage2_col105[11] <= fa_s1_c105_n515_s;
                    stage2_col105[12] <= fa_s1_c105_n516_s;
                    stage2_col105[13] <= fa_s1_c105_n517_s;
                    stage2_col105[14] <= stage1_col105[21];
                    stage2_col105[15] <= stage1_col105[22];
                    stage2_col106[0] <= fa_s1_c105_n511_c;
                    stage2_col106[1] <= fa_s1_c105_n512_c;
                    stage2_col106[2] <= fa_s1_c105_n513_c;
                    stage2_col106[3] <= fa_s1_c105_n514_c;
                    stage2_col106[4] <= fa_s1_c105_n515_c;
                    stage2_col106[5] <= fa_s1_c105_n516_c;
                    stage2_col106[6] <= fa_s1_c105_n517_c;
                    stage2_col106[7] <= fa_s1_c106_n518_s;
                    stage2_col106[8] <= fa_s1_c106_n519_s;
                    stage2_col106[9] <= fa_s1_c106_n520_s;
                    stage2_col106[10] <= fa_s1_c106_n521_s;
                    stage2_col106[11] <= fa_s1_c106_n522_s;
                    stage2_col106[12] <= fa_s1_c106_n523_s;
                    stage2_col106[13] <= fa_s1_c106_n524_s;
                    stage2_col107[0] <= fa_s1_c106_n518_c;
                    stage2_col107[1] <= fa_s1_c106_n519_c;
                    stage2_col107[2] <= fa_s1_c106_n520_c;
                    stage2_col107[3] <= fa_s1_c106_n521_c;
                    stage2_col107[4] <= fa_s1_c106_n522_c;
                    stage2_col107[5] <= fa_s1_c106_n523_c;
                    stage2_col107[6] <= fa_s1_c106_n524_c;
                    stage2_col107[7] <= fa_s1_c107_n525_s;
                    stage2_col107[8] <= fa_s1_c107_n526_s;
                    stage2_col107[9] <= fa_s1_c107_n527_s;
                    stage2_col107[10] <= fa_s1_c107_n528_s;
                    stage2_col107[11] <= fa_s1_c107_n529_s;
                    stage2_col107[12] <= fa_s1_c107_n530_s;
                    stage2_col107[13] <= fa_s1_c107_n531_s;
                    stage2_col107[14] <= stage1_col107[21];
                    stage2_col107[15] <= stage1_col107[22];
                    stage2_col108[0] <= fa_s1_c107_n525_c;
                    stage2_col108[1] <= fa_s1_c107_n526_c;
                    stage2_col108[2] <= fa_s1_c107_n527_c;
                    stage2_col108[3] <= fa_s1_c107_n528_c;
                    stage2_col108[4] <= fa_s1_c107_n529_c;
                    stage2_col108[5] <= fa_s1_c107_n530_c;
                    stage2_col108[6] <= fa_s1_c107_n531_c;
                    stage2_col108[7] <= fa_s1_c108_n532_s;
                    stage2_col108[8] <= fa_s1_c108_n533_s;
                    stage2_col108[9] <= fa_s1_c108_n534_s;
                    stage2_col108[10] <= fa_s1_c108_n535_s;
                    stage2_col108[11] <= fa_s1_c108_n536_s;
                    stage2_col108[12] <= fa_s1_c108_n537_s;
                    stage2_col108[13] <= fa_s1_c108_n538_s;
                    stage2_col109[0] <= fa_s1_c108_n532_c;
                    stage2_col109[1] <= fa_s1_c108_n533_c;
                    stage2_col109[2] <= fa_s1_c108_n534_c;
                    stage2_col109[3] <= fa_s1_c108_n535_c;
                    stage2_col109[4] <= fa_s1_c108_n536_c;
                    stage2_col109[5] <= fa_s1_c108_n537_c;
                    stage2_col109[6] <= fa_s1_c108_n538_c;
                    stage2_col109[7] <= fa_s1_c109_n539_s;
                    stage2_col109[8] <= fa_s1_c109_n540_s;
                    stage2_col109[9] <= fa_s1_c109_n541_s;
                    stage2_col109[10] <= fa_s1_c109_n542_s;
                    stage2_col109[11] <= fa_s1_c109_n543_s;
                    stage2_col109[12] <= fa_s1_c109_n544_s;
                    stage2_col109[13] <= fa_s1_c109_n545_s;
                    stage2_col109[14] <= stage1_col109[21];
                    stage2_col109[15] <= stage1_col109[22];
                    stage2_col110[0] <= fa_s1_c109_n539_c;
                    stage2_col110[1] <= fa_s1_c109_n540_c;
                    stage2_col110[2] <= fa_s1_c109_n541_c;
                    stage2_col110[3] <= fa_s1_c109_n542_c;
                    stage2_col110[4] <= fa_s1_c109_n543_c;
                    stage2_col110[5] <= fa_s1_c109_n544_c;
                    stage2_col110[6] <= fa_s1_c109_n545_c;
                    stage2_col110[7] <= fa_s1_c110_n546_s;
                    stage2_col110[8] <= fa_s1_c110_n547_s;
                    stage2_col110[9] <= fa_s1_c110_n548_s;
                    stage2_col110[10] <= fa_s1_c110_n549_s;
                    stage2_col110[11] <= fa_s1_c110_n550_s;
                    stage2_col110[12] <= fa_s1_c110_n551_s;
                    stage2_col110[13] <= fa_s1_c110_n552_s;
                    stage2_col111[0] <= fa_s1_c110_n546_c;
                    stage2_col111[1] <= fa_s1_c110_n547_c;
                    stage2_col111[2] <= fa_s1_c110_n548_c;
                    stage2_col111[3] <= fa_s1_c110_n549_c;
                    stage2_col111[4] <= fa_s1_c110_n550_c;
                    stage2_col111[5] <= fa_s1_c110_n551_c;
                    stage2_col111[6] <= fa_s1_c110_n552_c;
                    stage2_col111[7] <= fa_s1_c111_n553_s;
                    stage2_col111[8] <= fa_s1_c111_n554_s;
                    stage2_col111[9] <= fa_s1_c111_n555_s;
                    stage2_col111[10] <= fa_s1_c111_n556_s;
                    stage2_col111[11] <= fa_s1_c111_n557_s;
                    stage2_col111[12] <= fa_s1_c111_n558_s;
                    stage2_col111[13] <= fa_s1_c111_n559_s;
                    stage2_col111[14] <= stage1_col111[21];
                    stage2_col111[15] <= stage1_col111[22];
                    stage2_col112[0] <= fa_s1_c111_n553_c;
                    stage2_col112[1] <= fa_s1_c111_n554_c;
                    stage2_col112[2] <= fa_s1_c111_n555_c;
                    stage2_col112[3] <= fa_s1_c111_n556_c;
                    stage2_col112[4] <= fa_s1_c111_n557_c;
                    stage2_col112[5] <= fa_s1_c111_n558_c;
                    stage2_col112[6] <= fa_s1_c111_n559_c;
                    stage2_col112[7] <= fa_s1_c112_n560_s;
                    stage2_col112[8] <= fa_s1_c112_n561_s;
                    stage2_col112[9] <= fa_s1_c112_n562_s;
                    stage2_col112[10] <= fa_s1_c112_n563_s;
                    stage2_col112[11] <= fa_s1_c112_n564_s;
                    stage2_col112[12] <= fa_s1_c112_n565_s;
                    stage2_col112[13] <= fa_s1_c112_n566_s;
                    stage2_col113[0] <= fa_s1_c112_n560_c;
                    stage2_col113[1] <= fa_s1_c112_n561_c;
                    stage2_col113[2] <= fa_s1_c112_n562_c;
                    stage2_col113[3] <= fa_s1_c112_n563_c;
                    stage2_col113[4] <= fa_s1_c112_n564_c;
                    stage2_col113[5] <= fa_s1_c112_n565_c;
                    stage2_col113[6] <= fa_s1_c112_n566_c;
                    stage2_col113[7] <= fa_s1_c113_n567_s;
                    stage2_col113[8] <= fa_s1_c113_n568_s;
                    stage2_col113[9] <= fa_s1_c113_n569_s;
                    stage2_col113[10] <= fa_s1_c113_n570_s;
                    stage2_col113[11] <= fa_s1_c113_n571_s;
                    stage2_col113[12] <= fa_s1_c113_n572_s;
                    stage2_col113[13] <= fa_s1_c113_n573_s;
                    stage2_col113[14] <= stage1_col113[21];
                    stage2_col113[15] <= stage1_col113[22];
                    stage2_col114[0] <= fa_s1_c113_n567_c;
                    stage2_col114[1] <= fa_s1_c113_n568_c;
                    stage2_col114[2] <= fa_s1_c113_n569_c;
                    stage2_col114[3] <= fa_s1_c113_n570_c;
                    stage2_col114[4] <= fa_s1_c113_n571_c;
                    stage2_col114[5] <= fa_s1_c113_n572_c;
                    stage2_col114[6] <= fa_s1_c113_n573_c;
                    stage2_col114[7] <= fa_s1_c114_n574_s;
                    stage2_col114[8] <= fa_s1_c114_n575_s;
                    stage2_col114[9] <= fa_s1_c114_n576_s;
                    stage2_col114[10] <= fa_s1_c114_n577_s;
                    stage2_col114[11] <= fa_s1_c114_n578_s;
                    stage2_col114[12] <= fa_s1_c114_n579_s;
                    stage2_col114[13] <= fa_s1_c114_n580_s;
                    stage2_col115[0] <= fa_s1_c114_n574_c;
                    stage2_col115[1] <= fa_s1_c114_n575_c;
                    stage2_col115[2] <= fa_s1_c114_n576_c;
                    stage2_col115[3] <= fa_s1_c114_n577_c;
                    stage2_col115[4] <= fa_s1_c114_n578_c;
                    stage2_col115[5] <= fa_s1_c114_n579_c;
                    stage2_col115[6] <= fa_s1_c114_n580_c;
                    stage2_col115[7] <= fa_s1_c115_n581_s;
                    stage2_col115[8] <= fa_s1_c115_n582_s;
                    stage2_col115[9] <= fa_s1_c115_n583_s;
                    stage2_col115[10] <= fa_s1_c115_n584_s;
                    stage2_col115[11] <= fa_s1_c115_n585_s;
                    stage2_col115[12] <= fa_s1_c115_n586_s;
                    stage2_col115[13] <= fa_s1_c115_n587_s;
                    stage2_col115[14] <= stage1_col115[21];
                    stage2_col115[15] <= stage1_col115[22];
                    stage2_col116[0] <= fa_s1_c115_n581_c;
                    stage2_col116[1] <= fa_s1_c115_n582_c;
                    stage2_col116[2] <= fa_s1_c115_n583_c;
                    stage2_col116[3] <= fa_s1_c115_n584_c;
                    stage2_col116[4] <= fa_s1_c115_n585_c;
                    stage2_col116[5] <= fa_s1_c115_n586_c;
                    stage2_col116[6] <= fa_s1_c115_n587_c;
                    stage2_col116[7] <= fa_s1_c116_n588_s;
                    stage2_col116[8] <= fa_s1_c116_n589_s;
                    stage2_col116[9] <= fa_s1_c116_n590_s;
                    stage2_col116[10] <= fa_s1_c116_n591_s;
                    stage2_col116[11] <= fa_s1_c116_n592_s;
                    stage2_col116[12] <= fa_s1_c116_n593_s;
                    stage2_col116[13] <= fa_s1_c116_n594_s;
                    stage2_col117[0] <= fa_s1_c116_n588_c;
                    stage2_col117[1] <= fa_s1_c116_n589_c;
                    stage2_col117[2] <= fa_s1_c116_n590_c;
                    stage2_col117[3] <= fa_s1_c116_n591_c;
                    stage2_col117[4] <= fa_s1_c116_n592_c;
                    stage2_col117[5] <= fa_s1_c116_n593_c;
                    stage2_col117[6] <= fa_s1_c116_n594_c;
                    stage2_col117[7] <= fa_s1_c117_n595_s;
                    stage2_col117[8] <= fa_s1_c117_n596_s;
                    stage2_col117[9] <= fa_s1_c117_n597_s;
                    stage2_col117[10] <= fa_s1_c117_n598_s;
                    stage2_col117[11] <= fa_s1_c117_n599_s;
                    stage2_col117[12] <= fa_s1_c117_n600_s;
                    stage2_col117[13] <= fa_s1_c117_n601_s;
                    stage2_col117[14] <= stage1_col117[21];
                    stage2_col117[15] <= stage1_col117[22];
                    stage2_col118[0] <= fa_s1_c117_n595_c;
                    stage2_col118[1] <= fa_s1_c117_n596_c;
                    stage2_col118[2] <= fa_s1_c117_n597_c;
                    stage2_col118[3] <= fa_s1_c117_n598_c;
                    stage2_col118[4] <= fa_s1_c117_n599_c;
                    stage2_col118[5] <= fa_s1_c117_n600_c;
                    stage2_col118[6] <= fa_s1_c117_n601_c;
                    stage2_col118[7] <= fa_s1_c118_n602_s;
                    stage2_col118[8] <= fa_s1_c118_n603_s;
                    stage2_col118[9] <= fa_s1_c118_n604_s;
                    stage2_col118[10] <= fa_s1_c118_n605_s;
                    stage2_col118[11] <= fa_s1_c118_n606_s;
                    stage2_col118[12] <= fa_s1_c118_n607_s;
                    stage2_col118[13] <= fa_s1_c118_n608_s;
                    stage2_col119[0] <= fa_s1_c118_n602_c;
                    stage2_col119[1] <= fa_s1_c118_n603_c;
                    stage2_col119[2] <= fa_s1_c118_n604_c;
                    stage2_col119[3] <= fa_s1_c118_n605_c;
                    stage2_col119[4] <= fa_s1_c118_n606_c;
                    stage2_col119[5] <= fa_s1_c118_n607_c;
                    stage2_col119[6] <= fa_s1_c118_n608_c;
                    stage2_col119[7] <= fa_s1_c119_n609_s;
                    stage2_col119[8] <= fa_s1_c119_n610_s;
                    stage2_col119[9] <= fa_s1_c119_n611_s;
                    stage2_col119[10] <= fa_s1_c119_n612_s;
                    stage2_col119[11] <= fa_s1_c119_n613_s;
                    stage2_col119[12] <= fa_s1_c119_n614_s;
                    stage2_col119[13] <= fa_s1_c119_n615_s;
                    stage2_col119[14] <= stage1_col119[21];
                    stage2_col119[15] <= stage1_col119[22];
                    stage2_col120[0] <= fa_s1_c119_n609_c;
                    stage2_col120[1] <= fa_s1_c119_n610_c;
                    stage2_col120[2] <= fa_s1_c119_n611_c;
                    stage2_col120[3] <= fa_s1_c119_n612_c;
                    stage2_col120[4] <= fa_s1_c119_n613_c;
                    stage2_col120[5] <= fa_s1_c119_n614_c;
                    stage2_col120[6] <= fa_s1_c119_n615_c;
                    stage2_col120[7] <= fa_s1_c120_n616_s;
                    stage2_col120[8] <= fa_s1_c120_n617_s;
                    stage2_col120[9] <= fa_s1_c120_n618_s;
                    stage2_col120[10] <= fa_s1_c120_n619_s;
                    stage2_col120[11] <= fa_s1_c120_n620_s;
                    stage2_col120[12] <= fa_s1_c120_n621_s;
                    stage2_col120[13] <= fa_s1_c120_n622_s;
                    stage2_col121[0] <= fa_s1_c120_n616_c;
                    stage2_col121[1] <= fa_s1_c120_n617_c;
                    stage2_col121[2] <= fa_s1_c120_n618_c;
                    stage2_col121[3] <= fa_s1_c120_n619_c;
                    stage2_col121[4] <= fa_s1_c120_n620_c;
                    stage2_col121[5] <= fa_s1_c120_n621_c;
                    stage2_col121[6] <= fa_s1_c120_n622_c;
                    stage2_col121[7] <= fa_s1_c121_n623_s;
                    stage2_col121[8] <= fa_s1_c121_n624_s;
                    stage2_col121[9] <= fa_s1_c121_n625_s;
                    stage2_col121[10] <= fa_s1_c121_n626_s;
                    stage2_col121[11] <= fa_s1_c121_n627_s;
                    stage2_col121[12] <= fa_s1_c121_n628_s;
                    stage2_col121[13] <= fa_s1_c121_n629_s;
                    stage2_col121[14] <= stage1_col121[21];
                    stage2_col121[15] <= stage1_col121[22];
                    stage2_col122[0] <= fa_s1_c121_n623_c;
                    stage2_col122[1] <= fa_s1_c121_n624_c;
                    stage2_col122[2] <= fa_s1_c121_n625_c;
                    stage2_col122[3] <= fa_s1_c121_n626_c;
                    stage2_col122[4] <= fa_s1_c121_n627_c;
                    stage2_col122[5] <= fa_s1_c121_n628_c;
                    stage2_col122[6] <= fa_s1_c121_n629_c;
                    stage2_col122[7] <= fa_s1_c122_n630_s;
                    stage2_col122[8] <= fa_s1_c122_n631_s;
                    stage2_col122[9] <= fa_s1_c122_n632_s;
                    stage2_col122[10] <= fa_s1_c122_n633_s;
                    stage2_col122[11] <= fa_s1_c122_n634_s;
                    stage2_col122[12] <= fa_s1_c122_n635_s;
                    stage2_col122[13] <= fa_s1_c122_n636_s;
                    stage2_col123[0] <= fa_s1_c122_n630_c;
                    stage2_col123[1] <= fa_s1_c122_n631_c;
                    stage2_col123[2] <= fa_s1_c122_n632_c;
                    stage2_col123[3] <= fa_s1_c122_n633_c;
                    stage2_col123[4] <= fa_s1_c122_n634_c;
                    stage2_col123[5] <= fa_s1_c122_n635_c;
                    stage2_col123[6] <= fa_s1_c122_n636_c;
                    stage2_col123[7] <= fa_s1_c123_n637_s;
                    stage2_col123[8] <= fa_s1_c123_n638_s;
                    stage2_col123[9] <= fa_s1_c123_n639_s;
                    stage2_col123[10] <= fa_s1_c123_n640_s;
                    stage2_col123[11] <= fa_s1_c123_n641_s;
                    stage2_col123[12] <= fa_s1_c123_n642_s;
                    stage2_col123[13] <= fa_s1_c123_n643_s;
                    stage2_col123[14] <= stage1_col123[21];
                    stage2_col123[15] <= stage1_col123[22];
                    stage2_col124[0] <= fa_s1_c123_n637_c;
                    stage2_col124[1] <= fa_s1_c123_n638_c;
                    stage2_col124[2] <= fa_s1_c123_n639_c;
                    stage2_col124[3] <= fa_s1_c123_n640_c;
                    stage2_col124[4] <= fa_s1_c123_n641_c;
                    stage2_col124[5] <= fa_s1_c123_n642_c;
                    stage2_col124[6] <= fa_s1_c123_n643_c;
                    stage2_col124[7] <= fa_s1_c124_n644_s;
                    stage2_col124[8] <= fa_s1_c124_n645_s;
                    stage2_col124[9] <= fa_s1_c124_n646_s;
                    stage2_col124[10] <= fa_s1_c124_n647_s;
                    stage2_col124[11] <= fa_s1_c124_n648_s;
                    stage2_col124[12] <= fa_s1_c124_n649_s;
                    stage2_col124[13] <= fa_s1_c124_n650_s;
                    stage2_col125[0] <= fa_s1_c124_n644_c;
                    stage2_col125[1] <= fa_s1_c124_n645_c;
                    stage2_col125[2] <= fa_s1_c124_n646_c;
                    stage2_col125[3] <= fa_s1_c124_n647_c;
                    stage2_col125[4] <= fa_s1_c124_n648_c;
                    stage2_col125[5] <= fa_s1_c124_n649_c;
                    stage2_col125[6] <= fa_s1_c124_n650_c;
                    stage2_col125[7] <= fa_s1_c125_n651_s;
                    stage2_col125[8] <= fa_s1_c125_n652_s;
                    stage2_col125[9] <= fa_s1_c125_n653_s;
                    stage2_col125[10] <= fa_s1_c125_n654_s;
                    stage2_col125[11] <= fa_s1_c125_n655_s;
                    stage2_col125[12] <= fa_s1_c125_n656_s;
                    stage2_col125[13] <= fa_s1_c125_n657_s;
                    stage2_col125[14] <= stage1_col125[21];
                    stage2_col125[15] <= stage1_col125[22];
                    stage2_col126[0] <= fa_s1_c125_n651_c;
                    stage2_col126[1] <= fa_s1_c125_n652_c;
                    stage2_col126[2] <= fa_s1_c125_n653_c;
                    stage2_col126[3] <= fa_s1_c125_n654_c;
                    stage2_col126[4] <= fa_s1_c125_n655_c;
                    stage2_col126[5] <= fa_s1_c125_n656_c;
                    stage2_col126[6] <= fa_s1_c125_n657_c;
                    stage2_col126[7] <= fa_s1_c126_n658_s;
                    stage2_col126[8] <= fa_s1_c126_n659_s;
                    stage2_col126[9] <= fa_s1_c126_n660_s;
                    stage2_col126[10] <= fa_s1_c126_n661_s;
                    stage2_col126[11] <= fa_s1_c126_n662_s;
                    stage2_col126[12] <= fa_s1_c126_n663_s;
                    stage2_col126[13] <= fa_s1_c126_n664_s;
                    stage2_col127[0] <= fa_s1_c126_n658_c;
                    stage2_col127[1] <= fa_s1_c126_n659_c;
                    stage2_col127[2] <= fa_s1_c126_n660_c;
                    stage2_col127[3] <= fa_s1_c126_n661_c;
                    stage2_col127[4] <= fa_s1_c126_n662_c;
                    stage2_col127[5] <= fa_s1_c126_n663_c;
                    stage2_col127[6] <= fa_s1_c126_n664_c;
                    stage2_col127[7] <= stage1_col127[0];
                    stage2_col127[8] <= stage1_col127[1];
                    stage2_col127[9] <= stage1_col127[2];
                    stage2_col127[10] <= stage1_col127[3];
                    stage2_col127[11] <= stage1_col127[4];
                    stage2_col127[12] <= stage1_col127[5];
                    stage2_col127[13] <= stage1_col127[6];
                    stage2_col127[14] <= stage1_col127[7];
                    stage2_col127[15] <= stage1_col127[8];
                    stage2_col127[16] <= stage1_col127[9];
                    stage2_col127[17] <= stage1_col127[10];
                    stage2_col127[18] <= stage1_col127[11];
                    stage2_col127[19] <= stage1_col127[11];
                    stage2_col127[20] <= stage1_col127[11];
                    stage2_col127[21] <= stage1_col127[11];
                    stage2_col127[22] <= stage1_col127[11];
                    stage2_col127[23] <= stage1_col127[11];
                    stage2_col127[24] <= stage1_col127[11];
                    stage2_col127[25] <= stage1_col127[11];
                    stage2_col127[26] <= stage1_col127[11];
                    stage2_col127[27] <= stage1_col127[11];
                    stage2_col127[28] <= stage1_col127[11];
                    stage2_col127[29] <= stage1_col127[11];
                    stage2_col127[30] <= stage1_col127[11];
                    stage2_col127[31] <= stage1_col127[11];
                    stage2_col127[32] <= stage1_col127[11];
                    stage2_col127[33] <= stage1_col127[11];
                    stage2_col127[34] <= stage1_col127[11];
                    stage2_col127[35] <= stage1_col127[11];
                    stage2_col127[36] <= stage1_col127[11];
                    stage2_col127[37] <= stage1_col127[11];
                    stage2_col127[38] <= stage1_col127[11];
                    stage2_col127[39] <= stage1_col127[11];
                    stage2_col127[40] <= stage1_col127[11];
                    stage2_col127[41] <= stage1_col127[11];
                    stage2_col127[42] <= stage1_col127[11];
                    stage2_col127[43] <= stage1_col127[11];
                    stage2_col127[44] <= stage1_col127[11];
                    stage2_col127[45] <= stage1_col127[11];
                    stage2_col127[46] <= stage1_col127[11];
                    stage2_col127[47] <= stage1_col127[11];
                    stage2_col127[48] <= stage1_col127[11];
                    stage2_col127[49] <= stage1_col127[11];
                end
            end
        end else begin : gen_stage2_no_pipe
            // Combinational assignment
            always_comb begin
                stage2_col0[0] = stage1_col0[0];
                stage2_col1[0] = ha_s1_c1_n0_s;
                stage2_col2[0] = ha_s1_c1_n0_c;
                stage2_col2[1] = stage1_col2[0];
                stage2_col3[0] = fa_s1_c3_n0_s;
                stage2_col4[0] = fa_s1_c3_n0_c;
                stage2_col4[1] = stage1_col4[0];
                stage2_col4[2] = stage1_col4[1];
                stage2_col5[0] = stage1_col5[0];
                stage2_col5[1] = stage1_col5[1];
                stage2_col6[0] = fa_s1_c6_n1_s;
                stage2_col6[1] = stage1_col6[3];
                stage2_col7[0] = fa_s1_c6_n1_c;
                stage2_col7[1] = fa_s1_c7_n2_s;
                stage2_col8[0] = fa_s1_c7_n2_c;
                stage2_col8[1] = fa_s1_c8_n3_s;
                stage2_col9[0] = fa_s1_c8_n3_c;
                stage2_col9[1] = fa_s1_c9_n4_s;
                stage2_col9[2] = stage1_col9[3];
                stage2_col9[3] = stage1_col9[4];
                stage2_col10[0] = fa_s1_c9_n4_c;
                stage2_col10[1] = fa_s1_c10_n5_s;
                stage2_col10[2] = stage1_col10[3];
                stage2_col11[0] = fa_s1_c10_n5_c;
                stage2_col11[1] = fa_s1_c11_n6_s;
                stage2_col11[2] = stage1_col11[3];
                stage2_col12[0] = fa_s1_c11_n6_c;
                stage2_col12[1] = fa_s1_c12_n7_s;
                stage2_col12[2] = fa_s1_c12_n8_s;
                stage2_col13[0] = fa_s1_c12_n7_c;
                stage2_col13[1] = fa_s1_c12_n8_c;
                stage2_col13[2] = fa_s1_c13_n9_s;
                stage2_col13[3] = stage1_col13[3];
                stage2_col13[4] = stage1_col13[4];
                stage2_col14[0] = fa_s1_c13_n9_c;
                stage2_col14[1] = fa_s1_c14_n10_s;
                stage2_col14[2] = stage1_col14[3];
                stage2_col14[3] = stage1_col14[4];
                stage2_col15[0] = fa_s1_c14_n10_c;
                stage2_col15[1] = fa_s1_c15_n11_s;
                stage2_col15[2] = fa_s1_c15_n12_s;
                stage2_col15[3] = stage1_col15[6];
                stage2_col16[0] = fa_s1_c15_n11_c;
                stage2_col16[1] = fa_s1_c15_n12_c;
                stage2_col16[2] = fa_s1_c16_n13_s;
                stage2_col16[3] = fa_s1_c16_n14_s;
                stage2_col17[0] = fa_s1_c16_n13_c;
                stage2_col17[1] = fa_s1_c16_n14_c;
                stage2_col17[2] = fa_s1_c17_n15_s;
                stage2_col17[3] = fa_s1_c17_n16_s;
                stage2_col18[0] = fa_s1_c17_n15_c;
                stage2_col18[1] = fa_s1_c17_n16_c;
                stage2_col18[2] = fa_s1_c18_n17_s;
                stage2_col18[3] = fa_s1_c18_n18_s;
                stage2_col18[4] = stage1_col18[6];
                stage2_col18[5] = stage1_col18[7];
                stage2_col19[0] = fa_s1_c18_n17_c;
                stage2_col19[1] = fa_s1_c18_n18_c;
                stage2_col19[2] = fa_s1_c19_n19_s;
                stage2_col19[3] = fa_s1_c19_n20_s;
                stage2_col19[4] = stage1_col19[6];
                stage2_col20[0] = fa_s1_c19_n19_c;
                stage2_col20[1] = fa_s1_c19_n20_c;
                stage2_col20[2] = fa_s1_c20_n21_s;
                stage2_col20[3] = fa_s1_c20_n22_s;
                stage2_col20[4] = stage1_col20[6];
                stage2_col21[0] = fa_s1_c20_n21_c;
                stage2_col21[1] = fa_s1_c20_n22_c;
                stage2_col21[2] = fa_s1_c21_n23_s;
                stage2_col21[3] = fa_s1_c21_n24_s;
                stage2_col21[4] = fa_s1_c21_n25_s;
                stage2_col22[0] = fa_s1_c21_n23_c;
                stage2_col22[1] = fa_s1_c21_n24_c;
                stage2_col22[2] = fa_s1_c21_n25_c;
                stage2_col22[3] = fa_s1_c22_n26_s;
                stage2_col22[4] = fa_s1_c22_n27_s;
                stage2_col22[5] = stage1_col22[6];
                stage2_col22[6] = stage1_col22[7];
                stage2_col23[0] = fa_s1_c22_n26_c;
                stage2_col23[1] = fa_s1_c22_n27_c;
                stage2_col23[2] = fa_s1_c23_n28_s;
                stage2_col23[3] = fa_s1_c23_n29_s;
                stage2_col23[4] = stage1_col23[6];
                stage2_col23[5] = stage1_col23[7];
                stage2_col24[0] = fa_s1_c23_n28_c;
                stage2_col24[1] = fa_s1_c23_n29_c;
                stage2_col24[2] = fa_s1_c24_n30_s;
                stage2_col24[3] = fa_s1_c24_n31_s;
                stage2_col24[4] = fa_s1_c24_n32_s;
                stage2_col24[5] = stage1_col24[9];
                stage2_col25[0] = fa_s1_c24_n30_c;
                stage2_col25[1] = fa_s1_c24_n31_c;
                stage2_col25[2] = fa_s1_c24_n32_c;
                stage2_col25[3] = fa_s1_c25_n33_s;
                stage2_col25[4] = fa_s1_c25_n34_s;
                stage2_col25[5] = fa_s1_c25_n35_s;
                stage2_col26[0] = fa_s1_c25_n33_c;
                stage2_col26[1] = fa_s1_c25_n34_c;
                stage2_col26[2] = fa_s1_c25_n35_c;
                stage2_col26[3] = fa_s1_c26_n36_s;
                stage2_col26[4] = fa_s1_c26_n37_s;
                stage2_col26[5] = fa_s1_c26_n38_s;
                stage2_col27[0] = fa_s1_c26_n36_c;
                stage2_col27[1] = fa_s1_c26_n37_c;
                stage2_col27[2] = fa_s1_c26_n38_c;
                stage2_col27[3] = fa_s1_c27_n39_s;
                stage2_col27[4] = fa_s1_c27_n40_s;
                stage2_col27[5] = fa_s1_c27_n41_s;
                stage2_col27[6] = stage1_col27[9];
                stage2_col27[7] = stage1_col27[10];
                stage2_col28[0] = fa_s1_c27_n39_c;
                stage2_col28[1] = fa_s1_c27_n40_c;
                stage2_col28[2] = fa_s1_c27_n41_c;
                stage2_col28[3] = fa_s1_c28_n42_s;
                stage2_col28[4] = fa_s1_c28_n43_s;
                stage2_col28[5] = fa_s1_c28_n44_s;
                stage2_col28[6] = stage1_col28[9];
                stage2_col29[0] = fa_s1_c28_n42_c;
                stage2_col29[1] = fa_s1_c28_n43_c;
                stage2_col29[2] = fa_s1_c28_n44_c;
                stage2_col29[3] = fa_s1_c29_n45_s;
                stage2_col29[4] = fa_s1_c29_n46_s;
                stage2_col29[5] = fa_s1_c29_n47_s;
                stage2_col29[6] = stage1_col29[9];
                stage2_col30[0] = fa_s1_c29_n45_c;
                stage2_col30[1] = fa_s1_c29_n46_c;
                stage2_col30[2] = fa_s1_c29_n47_c;
                stage2_col30[3] = fa_s1_c30_n48_s;
                stage2_col30[4] = fa_s1_c30_n49_s;
                stage2_col30[5] = fa_s1_c30_n50_s;
                stage2_col30[6] = fa_s1_c30_n51_s;
                stage2_col31[0] = fa_s1_c30_n48_c;
                stage2_col31[1] = fa_s1_c30_n49_c;
                stage2_col31[2] = fa_s1_c30_n50_c;
                stage2_col31[3] = fa_s1_c30_n51_c;
                stage2_col31[4] = fa_s1_c31_n52_s;
                stage2_col31[5] = fa_s1_c31_n53_s;
                stage2_col31[6] = fa_s1_c31_n54_s;
                stage2_col31[7] = stage1_col31[9];
                stage2_col31[8] = stage1_col31[10];
                stage2_col32[0] = fa_s1_c31_n52_c;
                stage2_col32[1] = fa_s1_c31_n53_c;
                stage2_col32[2] = fa_s1_c31_n54_c;
                stage2_col32[3] = fa_s1_c32_n55_s;
                stage2_col32[4] = fa_s1_c32_n56_s;
                stage2_col32[5] = fa_s1_c32_n57_s;
                stage2_col32[6] = stage1_col32[9];
                stage2_col32[7] = stage1_col32[10];
                stage2_col33[0] = fa_s1_c32_n55_c;
                stage2_col33[1] = fa_s1_c32_n56_c;
                stage2_col33[2] = fa_s1_c32_n57_c;
                stage2_col33[3] = fa_s1_c33_n58_s;
                stage2_col33[4] = fa_s1_c33_n59_s;
                stage2_col33[5] = fa_s1_c33_n60_s;
                stage2_col33[6] = fa_s1_c33_n61_s;
                stage2_col33[7] = stage1_col33[12];
                stage2_col34[0] = fa_s1_c33_n58_c;
                stage2_col34[1] = fa_s1_c33_n59_c;
                stage2_col34[2] = fa_s1_c33_n60_c;
                stage2_col34[3] = fa_s1_c33_n61_c;
                stage2_col34[4] = fa_s1_c34_n62_s;
                stage2_col34[5] = fa_s1_c34_n63_s;
                stage2_col34[6] = fa_s1_c34_n64_s;
                stage2_col34[7] = fa_s1_c34_n65_s;
                stage2_col35[0] = fa_s1_c34_n62_c;
                stage2_col35[1] = fa_s1_c34_n63_c;
                stage2_col35[2] = fa_s1_c34_n64_c;
                stage2_col35[3] = fa_s1_c34_n65_c;
                stage2_col35[4] = fa_s1_c35_n66_s;
                stage2_col35[5] = fa_s1_c35_n67_s;
                stage2_col35[6] = fa_s1_c35_n68_s;
                stage2_col35[7] = fa_s1_c35_n69_s;
                stage2_col36[0] = fa_s1_c35_n66_c;
                stage2_col36[1] = fa_s1_c35_n67_c;
                stage2_col36[2] = fa_s1_c35_n68_c;
                stage2_col36[3] = fa_s1_c35_n69_c;
                stage2_col36[4] = fa_s1_c36_n70_s;
                stage2_col36[5] = fa_s1_c36_n71_s;
                stage2_col36[6] = fa_s1_c36_n72_s;
                stage2_col36[7] = fa_s1_c36_n73_s;
                stage2_col36[8] = stage1_col36[12];
                stage2_col36[9] = stage1_col36[13];
                stage2_col37[0] = fa_s1_c36_n70_c;
                stage2_col37[1] = fa_s1_c36_n71_c;
                stage2_col37[2] = fa_s1_c36_n72_c;
                stage2_col37[3] = fa_s1_c36_n73_c;
                stage2_col37[4] = fa_s1_c37_n74_s;
                stage2_col37[5] = fa_s1_c37_n75_s;
                stage2_col37[6] = fa_s1_c37_n76_s;
                stage2_col37[7] = fa_s1_c37_n77_s;
                stage2_col37[8] = stage1_col37[12];
                stage2_col38[0] = fa_s1_c37_n74_c;
                stage2_col38[1] = fa_s1_c37_n75_c;
                stage2_col38[2] = fa_s1_c37_n76_c;
                stage2_col38[3] = fa_s1_c37_n77_c;
                stage2_col38[4] = fa_s1_c38_n78_s;
                stage2_col38[5] = fa_s1_c38_n79_s;
                stage2_col38[6] = fa_s1_c38_n80_s;
                stage2_col38[7] = fa_s1_c38_n81_s;
                stage2_col38[8] = stage1_col38[12];
                stage2_col39[0] = fa_s1_c38_n78_c;
                stage2_col39[1] = fa_s1_c38_n79_c;
                stage2_col39[2] = fa_s1_c38_n80_c;
                stage2_col39[3] = fa_s1_c38_n81_c;
                stage2_col39[4] = fa_s1_c39_n82_s;
                stage2_col39[5] = fa_s1_c39_n83_s;
                stage2_col39[6] = fa_s1_c39_n84_s;
                stage2_col39[7] = fa_s1_c39_n85_s;
                stage2_col39[8] = fa_s1_c39_n86_s;
                stage2_col40[0] = fa_s1_c39_n82_c;
                stage2_col40[1] = fa_s1_c39_n83_c;
                stage2_col40[2] = fa_s1_c39_n84_c;
                stage2_col40[3] = fa_s1_c39_n85_c;
                stage2_col40[4] = fa_s1_c39_n86_c;
                stage2_col40[5] = fa_s1_c40_n87_s;
                stage2_col40[6] = fa_s1_c40_n88_s;
                stage2_col40[7] = fa_s1_c40_n89_s;
                stage2_col40[8] = fa_s1_c40_n90_s;
                stage2_col40[9] = stage1_col40[12];
                stage2_col40[10] = stage1_col40[13];
                stage2_col41[0] = fa_s1_c40_n87_c;
                stage2_col41[1] = fa_s1_c40_n88_c;
                stage2_col41[2] = fa_s1_c40_n89_c;
                stage2_col41[3] = fa_s1_c40_n90_c;
                stage2_col41[4] = fa_s1_c41_n91_s;
                stage2_col41[5] = fa_s1_c41_n92_s;
                stage2_col41[6] = fa_s1_c41_n93_s;
                stage2_col41[7] = fa_s1_c41_n94_s;
                stage2_col41[8] = stage1_col41[12];
                stage2_col41[9] = stage1_col41[13];
                stage2_col42[0] = fa_s1_c41_n91_c;
                stage2_col42[1] = fa_s1_c41_n92_c;
                stage2_col42[2] = fa_s1_c41_n93_c;
                stage2_col42[3] = fa_s1_c41_n94_c;
                stage2_col42[4] = fa_s1_c42_n95_s;
                stage2_col42[5] = fa_s1_c42_n96_s;
                stage2_col42[6] = fa_s1_c42_n97_s;
                stage2_col42[7] = fa_s1_c42_n98_s;
                stage2_col42[8] = fa_s1_c42_n99_s;
                stage2_col42[9] = stage1_col42[15];
                stage2_col43[0] = fa_s1_c42_n95_c;
                stage2_col43[1] = fa_s1_c42_n96_c;
                stage2_col43[2] = fa_s1_c42_n97_c;
                stage2_col43[3] = fa_s1_c42_n98_c;
                stage2_col43[4] = fa_s1_c42_n99_c;
                stage2_col43[5] = fa_s1_c43_n100_s;
                stage2_col43[6] = fa_s1_c43_n101_s;
                stage2_col43[7] = fa_s1_c43_n102_s;
                stage2_col43[8] = fa_s1_c43_n103_s;
                stage2_col43[9] = fa_s1_c43_n104_s;
                stage2_col44[0] = fa_s1_c43_n100_c;
                stage2_col44[1] = fa_s1_c43_n101_c;
                stage2_col44[2] = fa_s1_c43_n102_c;
                stage2_col44[3] = fa_s1_c43_n103_c;
                stage2_col44[4] = fa_s1_c43_n104_c;
                stage2_col44[5] = fa_s1_c44_n105_s;
                stage2_col44[6] = fa_s1_c44_n106_s;
                stage2_col44[7] = fa_s1_c44_n107_s;
                stage2_col44[8] = fa_s1_c44_n108_s;
                stage2_col44[9] = fa_s1_c44_n109_s;
                stage2_col45[0] = fa_s1_c44_n105_c;
                stage2_col45[1] = fa_s1_c44_n106_c;
                stage2_col45[2] = fa_s1_c44_n107_c;
                stage2_col45[3] = fa_s1_c44_n108_c;
                stage2_col45[4] = fa_s1_c44_n109_c;
                stage2_col45[5] = fa_s1_c45_n110_s;
                stage2_col45[6] = fa_s1_c45_n111_s;
                stage2_col45[7] = fa_s1_c45_n112_s;
                stage2_col45[8] = fa_s1_c45_n113_s;
                stage2_col45[9] = fa_s1_c45_n114_s;
                stage2_col45[10] = stage1_col45[15];
                stage2_col45[11] = stage1_col45[16];
                stage2_col46[0] = fa_s1_c45_n110_c;
                stage2_col46[1] = fa_s1_c45_n111_c;
                stage2_col46[2] = fa_s1_c45_n112_c;
                stage2_col46[3] = fa_s1_c45_n113_c;
                stage2_col46[4] = fa_s1_c45_n114_c;
                stage2_col46[5] = fa_s1_c46_n115_s;
                stage2_col46[6] = fa_s1_c46_n116_s;
                stage2_col46[7] = fa_s1_c46_n117_s;
                stage2_col46[8] = fa_s1_c46_n118_s;
                stage2_col46[9] = fa_s1_c46_n119_s;
                stage2_col46[10] = stage1_col46[15];
                stage2_col47[0] = fa_s1_c46_n115_c;
                stage2_col47[1] = fa_s1_c46_n116_c;
                stage2_col47[2] = fa_s1_c46_n117_c;
                stage2_col47[3] = fa_s1_c46_n118_c;
                stage2_col47[4] = fa_s1_c46_n119_c;
                stage2_col47[5] = fa_s1_c47_n120_s;
                stage2_col47[6] = fa_s1_c47_n121_s;
                stage2_col47[7] = fa_s1_c47_n122_s;
                stage2_col47[8] = fa_s1_c47_n123_s;
                stage2_col47[9] = fa_s1_c47_n124_s;
                stage2_col47[10] = stage1_col47[15];
                stage2_col48[0] = fa_s1_c47_n120_c;
                stage2_col48[1] = fa_s1_c47_n121_c;
                stage2_col48[2] = fa_s1_c47_n122_c;
                stage2_col48[3] = fa_s1_c47_n123_c;
                stage2_col48[4] = fa_s1_c47_n124_c;
                stage2_col48[5] = fa_s1_c48_n125_s;
                stage2_col48[6] = fa_s1_c48_n126_s;
                stage2_col48[7] = fa_s1_c48_n127_s;
                stage2_col48[8] = fa_s1_c48_n128_s;
                stage2_col48[9] = fa_s1_c48_n129_s;
                stage2_col48[10] = fa_s1_c48_n130_s;
                stage2_col49[0] = fa_s1_c48_n125_c;
                stage2_col49[1] = fa_s1_c48_n126_c;
                stage2_col49[2] = fa_s1_c48_n127_c;
                stage2_col49[3] = fa_s1_c48_n128_c;
                stage2_col49[4] = fa_s1_c48_n129_c;
                stage2_col49[5] = fa_s1_c48_n130_c;
                stage2_col49[6] = fa_s1_c49_n131_s;
                stage2_col49[7] = fa_s1_c49_n132_s;
                stage2_col49[8] = fa_s1_c49_n133_s;
                stage2_col49[9] = fa_s1_c49_n134_s;
                stage2_col49[10] = fa_s1_c49_n135_s;
                stage2_col49[11] = stage1_col49[15];
                stage2_col49[12] = stage1_col49[16];
                stage2_col50[0] = fa_s1_c49_n131_c;
                stage2_col50[1] = fa_s1_c49_n132_c;
                stage2_col50[2] = fa_s1_c49_n133_c;
                stage2_col50[3] = fa_s1_c49_n134_c;
                stage2_col50[4] = fa_s1_c49_n135_c;
                stage2_col50[5] = fa_s1_c50_n136_s;
                stage2_col50[6] = fa_s1_c50_n137_s;
                stage2_col50[7] = fa_s1_c50_n138_s;
                stage2_col50[8] = fa_s1_c50_n139_s;
                stage2_col50[9] = fa_s1_c50_n140_s;
                stage2_col50[10] = stage1_col50[15];
                stage2_col50[11] = stage1_col50[16];
                stage2_col51[0] = fa_s1_c50_n136_c;
                stage2_col51[1] = fa_s1_c50_n137_c;
                stage2_col51[2] = fa_s1_c50_n138_c;
                stage2_col51[3] = fa_s1_c50_n139_c;
                stage2_col51[4] = fa_s1_c50_n140_c;
                stage2_col51[5] = fa_s1_c51_n141_s;
                stage2_col51[6] = fa_s1_c51_n142_s;
                stage2_col51[7] = fa_s1_c51_n143_s;
                stage2_col51[8] = fa_s1_c51_n144_s;
                stage2_col51[9] = fa_s1_c51_n145_s;
                stage2_col51[10] = fa_s1_c51_n146_s;
                stage2_col51[11] = stage1_col51[18];
                stage2_col52[0] = fa_s1_c51_n141_c;
                stage2_col52[1] = fa_s1_c51_n142_c;
                stage2_col52[2] = fa_s1_c51_n143_c;
                stage2_col52[3] = fa_s1_c51_n144_c;
                stage2_col52[4] = fa_s1_c51_n145_c;
                stage2_col52[5] = fa_s1_c51_n146_c;
                stage2_col52[6] = fa_s1_c52_n147_s;
                stage2_col52[7] = fa_s1_c52_n148_s;
                stage2_col52[8] = fa_s1_c52_n149_s;
                stage2_col52[9] = fa_s1_c52_n150_s;
                stage2_col52[10] = fa_s1_c52_n151_s;
                stage2_col52[11] = fa_s1_c52_n152_s;
                stage2_col53[0] = fa_s1_c52_n147_c;
                stage2_col53[1] = fa_s1_c52_n148_c;
                stage2_col53[2] = fa_s1_c52_n149_c;
                stage2_col53[3] = fa_s1_c52_n150_c;
                stage2_col53[4] = fa_s1_c52_n151_c;
                stage2_col53[5] = fa_s1_c52_n152_c;
                stage2_col53[6] = fa_s1_c53_n153_s;
                stage2_col53[7] = fa_s1_c53_n154_s;
                stage2_col53[8] = fa_s1_c53_n155_s;
                stage2_col53[9] = fa_s1_c53_n156_s;
                stage2_col53[10] = fa_s1_c53_n157_s;
                stage2_col53[11] = fa_s1_c53_n158_s;
                stage2_col54[0] = fa_s1_c53_n153_c;
                stage2_col54[1] = fa_s1_c53_n154_c;
                stage2_col54[2] = fa_s1_c53_n155_c;
                stage2_col54[3] = fa_s1_c53_n156_c;
                stage2_col54[4] = fa_s1_c53_n157_c;
                stage2_col54[5] = fa_s1_c53_n158_c;
                stage2_col54[6] = fa_s1_c54_n159_s;
                stage2_col54[7] = fa_s1_c54_n160_s;
                stage2_col54[8] = fa_s1_c54_n161_s;
                stage2_col54[9] = fa_s1_c54_n162_s;
                stage2_col54[10] = fa_s1_c54_n163_s;
                stage2_col54[11] = fa_s1_c54_n164_s;
                stage2_col54[12] = stage1_col54[18];
                stage2_col54[13] = stage1_col54[19];
                stage2_col55[0] = fa_s1_c54_n159_c;
                stage2_col55[1] = fa_s1_c54_n160_c;
                stage2_col55[2] = fa_s1_c54_n161_c;
                stage2_col55[3] = fa_s1_c54_n162_c;
                stage2_col55[4] = fa_s1_c54_n163_c;
                stage2_col55[5] = fa_s1_c54_n164_c;
                stage2_col55[6] = fa_s1_c55_n165_s;
                stage2_col55[7] = fa_s1_c55_n166_s;
                stage2_col55[8] = fa_s1_c55_n167_s;
                stage2_col55[9] = fa_s1_c55_n168_s;
                stage2_col55[10] = fa_s1_c55_n169_s;
                stage2_col55[11] = fa_s1_c55_n170_s;
                stage2_col55[12] = stage1_col55[18];
                stage2_col56[0] = fa_s1_c55_n165_c;
                stage2_col56[1] = fa_s1_c55_n166_c;
                stage2_col56[2] = fa_s1_c55_n167_c;
                stage2_col56[3] = fa_s1_c55_n168_c;
                stage2_col56[4] = fa_s1_c55_n169_c;
                stage2_col56[5] = fa_s1_c55_n170_c;
                stage2_col56[6] = fa_s1_c56_n171_s;
                stage2_col56[7] = fa_s1_c56_n172_s;
                stage2_col56[8] = fa_s1_c56_n173_s;
                stage2_col56[9] = fa_s1_c56_n174_s;
                stage2_col56[10] = fa_s1_c56_n175_s;
                stage2_col56[11] = fa_s1_c56_n176_s;
                stage2_col56[12] = stage1_col56[18];
                stage2_col57[0] = fa_s1_c56_n171_c;
                stage2_col57[1] = fa_s1_c56_n172_c;
                stage2_col57[2] = fa_s1_c56_n173_c;
                stage2_col57[3] = fa_s1_c56_n174_c;
                stage2_col57[4] = fa_s1_c56_n175_c;
                stage2_col57[5] = fa_s1_c56_n176_c;
                stage2_col57[6] = fa_s1_c57_n177_s;
                stage2_col57[7] = fa_s1_c57_n178_s;
                stage2_col57[8] = fa_s1_c57_n179_s;
                stage2_col57[9] = fa_s1_c57_n180_s;
                stage2_col57[10] = fa_s1_c57_n181_s;
                stage2_col57[11] = fa_s1_c57_n182_s;
                stage2_col57[12] = fa_s1_c57_n183_s;
                stage2_col58[0] = fa_s1_c57_n177_c;
                stage2_col58[1] = fa_s1_c57_n178_c;
                stage2_col58[2] = fa_s1_c57_n179_c;
                stage2_col58[3] = fa_s1_c57_n180_c;
                stage2_col58[4] = fa_s1_c57_n181_c;
                stage2_col58[5] = fa_s1_c57_n182_c;
                stage2_col58[6] = fa_s1_c57_n183_c;
                stage2_col58[7] = fa_s1_c58_n184_s;
                stage2_col58[8] = fa_s1_c58_n185_s;
                stage2_col58[9] = fa_s1_c58_n186_s;
                stage2_col58[10] = fa_s1_c58_n187_s;
                stage2_col58[11] = fa_s1_c58_n188_s;
                stage2_col58[12] = fa_s1_c58_n189_s;
                stage2_col58[13] = stage1_col58[18];
                stage2_col58[14] = stage1_col58[19];
                stage2_col59[0] = fa_s1_c58_n184_c;
                stage2_col59[1] = fa_s1_c58_n185_c;
                stage2_col59[2] = fa_s1_c58_n186_c;
                stage2_col59[3] = fa_s1_c58_n187_c;
                stage2_col59[4] = fa_s1_c58_n188_c;
                stage2_col59[5] = fa_s1_c58_n189_c;
                stage2_col59[6] = fa_s1_c59_n190_s;
                stage2_col59[7] = fa_s1_c59_n191_s;
                stage2_col59[8] = fa_s1_c59_n192_s;
                stage2_col59[9] = fa_s1_c59_n193_s;
                stage2_col59[10] = fa_s1_c59_n194_s;
                stage2_col59[11] = fa_s1_c59_n195_s;
                stage2_col59[12] = stage1_col59[18];
                stage2_col59[13] = stage1_col59[19];
                stage2_col60[0] = fa_s1_c59_n190_c;
                stage2_col60[1] = fa_s1_c59_n191_c;
                stage2_col60[2] = fa_s1_c59_n192_c;
                stage2_col60[3] = fa_s1_c59_n193_c;
                stage2_col60[4] = fa_s1_c59_n194_c;
                stage2_col60[5] = fa_s1_c59_n195_c;
                stage2_col60[6] = fa_s1_c60_n196_s;
                stage2_col60[7] = fa_s1_c60_n197_s;
                stage2_col60[8] = fa_s1_c60_n198_s;
                stage2_col60[9] = fa_s1_c60_n199_s;
                stage2_col60[10] = fa_s1_c60_n200_s;
                stage2_col60[11] = fa_s1_c60_n201_s;
                stage2_col60[12] = fa_s1_c60_n202_s;
                stage2_col60[13] = stage1_col60[21];
                stage2_col61[0] = fa_s1_c60_n196_c;
                stage2_col61[1] = fa_s1_c60_n197_c;
                stage2_col61[2] = fa_s1_c60_n198_c;
                stage2_col61[3] = fa_s1_c60_n199_c;
                stage2_col61[4] = fa_s1_c60_n200_c;
                stage2_col61[5] = fa_s1_c60_n201_c;
                stage2_col61[6] = fa_s1_c60_n202_c;
                stage2_col61[7] = fa_s1_c61_n203_s;
                stage2_col61[8] = fa_s1_c61_n204_s;
                stage2_col61[9] = fa_s1_c61_n205_s;
                stage2_col61[10] = fa_s1_c61_n206_s;
                stage2_col61[11] = fa_s1_c61_n207_s;
                stage2_col61[12] = fa_s1_c61_n208_s;
                stage2_col61[13] = fa_s1_c61_n209_s;
                stage2_col62[0] = fa_s1_c61_n203_c;
                stage2_col62[1] = fa_s1_c61_n204_c;
                stage2_col62[2] = fa_s1_c61_n205_c;
                stage2_col62[3] = fa_s1_c61_n206_c;
                stage2_col62[4] = fa_s1_c61_n207_c;
                stage2_col62[5] = fa_s1_c61_n208_c;
                stage2_col62[6] = fa_s1_c61_n209_c;
                stage2_col62[7] = fa_s1_c62_n210_s;
                stage2_col62[8] = fa_s1_c62_n211_s;
                stage2_col62[9] = fa_s1_c62_n212_s;
                stage2_col62[10] = fa_s1_c62_n213_s;
                stage2_col62[11] = fa_s1_c62_n214_s;
                stage2_col62[12] = fa_s1_c62_n215_s;
                stage2_col62[13] = fa_s1_c62_n216_s;
                stage2_col63[0] = fa_s1_c62_n210_c;
                stage2_col63[1] = fa_s1_c62_n211_c;
                stage2_col63[2] = fa_s1_c62_n212_c;
                stage2_col63[3] = fa_s1_c62_n213_c;
                stage2_col63[4] = fa_s1_c62_n214_c;
                stage2_col63[5] = fa_s1_c62_n215_c;
                stage2_col63[6] = fa_s1_c62_n216_c;
                stage2_col63[7] = fa_s1_c63_n217_s;
                stage2_col63[8] = fa_s1_c63_n218_s;
                stage2_col63[9] = fa_s1_c63_n219_s;
                stage2_col63[10] = fa_s1_c63_n220_s;
                stage2_col63[11] = fa_s1_c63_n221_s;
                stage2_col63[12] = fa_s1_c63_n222_s;
                stage2_col63[13] = fa_s1_c63_n223_s;
                stage2_col63[14] = stage1_col63[21];
                stage2_col63[15] = stage1_col63[22];
                stage2_col64[0] = fa_s1_c63_n217_c;
                stage2_col64[1] = fa_s1_c63_n218_c;
                stage2_col64[2] = fa_s1_c63_n219_c;
                stage2_col64[3] = fa_s1_c63_n220_c;
                stage2_col64[4] = fa_s1_c63_n221_c;
                stage2_col64[5] = fa_s1_c63_n222_c;
                stage2_col64[6] = fa_s1_c63_n223_c;
                stage2_col64[7] = fa_s1_c64_n224_s;
                stage2_col64[8] = fa_s1_c64_n225_s;
                stage2_col64[9] = fa_s1_c64_n226_s;
                stage2_col64[10] = fa_s1_c64_n227_s;
                stage2_col64[11] = fa_s1_c64_n228_s;
                stage2_col64[12] = fa_s1_c64_n229_s;
                stage2_col64[13] = fa_s1_c64_n230_s;
                stage2_col65[0] = fa_s1_c64_n224_c;
                stage2_col65[1] = fa_s1_c64_n225_c;
                stage2_col65[2] = fa_s1_c64_n226_c;
                stage2_col65[3] = fa_s1_c64_n227_c;
                stage2_col65[4] = fa_s1_c64_n228_c;
                stage2_col65[5] = fa_s1_c64_n229_c;
                stage2_col65[6] = fa_s1_c64_n230_c;
                stage2_col65[7] = fa_s1_c65_n231_s;
                stage2_col65[8] = fa_s1_c65_n232_s;
                stage2_col65[9] = fa_s1_c65_n233_s;
                stage2_col65[10] = fa_s1_c65_n234_s;
                stage2_col65[11] = fa_s1_c65_n235_s;
                stage2_col65[12] = fa_s1_c65_n236_s;
                stage2_col65[13] = fa_s1_c65_n237_s;
                stage2_col65[14] = stage1_col65[21];
                stage2_col65[15] = stage1_col65[22];
                stage2_col66[0] = fa_s1_c65_n231_c;
                stage2_col66[1] = fa_s1_c65_n232_c;
                stage2_col66[2] = fa_s1_c65_n233_c;
                stage2_col66[3] = fa_s1_c65_n234_c;
                stage2_col66[4] = fa_s1_c65_n235_c;
                stage2_col66[5] = fa_s1_c65_n236_c;
                stage2_col66[6] = fa_s1_c65_n237_c;
                stage2_col66[7] = fa_s1_c66_n238_s;
                stage2_col66[8] = fa_s1_c66_n239_s;
                stage2_col66[9] = fa_s1_c66_n240_s;
                stage2_col66[10] = fa_s1_c66_n241_s;
                stage2_col66[11] = fa_s1_c66_n242_s;
                stage2_col66[12] = fa_s1_c66_n243_s;
                stage2_col66[13] = fa_s1_c66_n244_s;
                stage2_col67[0] = fa_s1_c66_n238_c;
                stage2_col67[1] = fa_s1_c66_n239_c;
                stage2_col67[2] = fa_s1_c66_n240_c;
                stage2_col67[3] = fa_s1_c66_n241_c;
                stage2_col67[4] = fa_s1_c66_n242_c;
                stage2_col67[5] = fa_s1_c66_n243_c;
                stage2_col67[6] = fa_s1_c66_n244_c;
                stage2_col67[7] = fa_s1_c67_n245_s;
                stage2_col67[8] = fa_s1_c67_n246_s;
                stage2_col67[9] = fa_s1_c67_n247_s;
                stage2_col67[10] = fa_s1_c67_n248_s;
                stage2_col67[11] = fa_s1_c67_n249_s;
                stage2_col67[12] = fa_s1_c67_n250_s;
                stage2_col67[13] = fa_s1_c67_n251_s;
                stage2_col67[14] = stage1_col67[21];
                stage2_col67[15] = stage1_col67[22];
                stage2_col68[0] = fa_s1_c67_n245_c;
                stage2_col68[1] = fa_s1_c67_n246_c;
                stage2_col68[2] = fa_s1_c67_n247_c;
                stage2_col68[3] = fa_s1_c67_n248_c;
                stage2_col68[4] = fa_s1_c67_n249_c;
                stage2_col68[5] = fa_s1_c67_n250_c;
                stage2_col68[6] = fa_s1_c67_n251_c;
                stage2_col68[7] = fa_s1_c68_n252_s;
                stage2_col68[8] = fa_s1_c68_n253_s;
                stage2_col68[9] = fa_s1_c68_n254_s;
                stage2_col68[10] = fa_s1_c68_n255_s;
                stage2_col68[11] = fa_s1_c68_n256_s;
                stage2_col68[12] = fa_s1_c68_n257_s;
                stage2_col68[13] = fa_s1_c68_n258_s;
                stage2_col69[0] = fa_s1_c68_n252_c;
                stage2_col69[1] = fa_s1_c68_n253_c;
                stage2_col69[2] = fa_s1_c68_n254_c;
                stage2_col69[3] = fa_s1_c68_n255_c;
                stage2_col69[4] = fa_s1_c68_n256_c;
                stage2_col69[5] = fa_s1_c68_n257_c;
                stage2_col69[6] = fa_s1_c68_n258_c;
                stage2_col69[7] = fa_s1_c69_n259_s;
                stage2_col69[8] = fa_s1_c69_n260_s;
                stage2_col69[9] = fa_s1_c69_n261_s;
                stage2_col69[10] = fa_s1_c69_n262_s;
                stage2_col69[11] = fa_s1_c69_n263_s;
                stage2_col69[12] = fa_s1_c69_n264_s;
                stage2_col69[13] = fa_s1_c69_n265_s;
                stage2_col69[14] = stage1_col69[21];
                stage2_col69[15] = stage1_col69[22];
                stage2_col70[0] = fa_s1_c69_n259_c;
                stage2_col70[1] = fa_s1_c69_n260_c;
                stage2_col70[2] = fa_s1_c69_n261_c;
                stage2_col70[3] = fa_s1_c69_n262_c;
                stage2_col70[4] = fa_s1_c69_n263_c;
                stage2_col70[5] = fa_s1_c69_n264_c;
                stage2_col70[6] = fa_s1_c69_n265_c;
                stage2_col70[7] = fa_s1_c70_n266_s;
                stage2_col70[8] = fa_s1_c70_n267_s;
                stage2_col70[9] = fa_s1_c70_n268_s;
                stage2_col70[10] = fa_s1_c70_n269_s;
                stage2_col70[11] = fa_s1_c70_n270_s;
                stage2_col70[12] = fa_s1_c70_n271_s;
                stage2_col70[13] = fa_s1_c70_n272_s;
                stage2_col71[0] = fa_s1_c70_n266_c;
                stage2_col71[1] = fa_s1_c70_n267_c;
                stage2_col71[2] = fa_s1_c70_n268_c;
                stage2_col71[3] = fa_s1_c70_n269_c;
                stage2_col71[4] = fa_s1_c70_n270_c;
                stage2_col71[5] = fa_s1_c70_n271_c;
                stage2_col71[6] = fa_s1_c70_n272_c;
                stage2_col71[7] = fa_s1_c71_n273_s;
                stage2_col71[8] = fa_s1_c71_n274_s;
                stage2_col71[9] = fa_s1_c71_n275_s;
                stage2_col71[10] = fa_s1_c71_n276_s;
                stage2_col71[11] = fa_s1_c71_n277_s;
                stage2_col71[12] = fa_s1_c71_n278_s;
                stage2_col71[13] = fa_s1_c71_n279_s;
                stage2_col71[14] = stage1_col71[21];
                stage2_col71[15] = stage1_col71[22];
                stage2_col72[0] = fa_s1_c71_n273_c;
                stage2_col72[1] = fa_s1_c71_n274_c;
                stage2_col72[2] = fa_s1_c71_n275_c;
                stage2_col72[3] = fa_s1_c71_n276_c;
                stage2_col72[4] = fa_s1_c71_n277_c;
                stage2_col72[5] = fa_s1_c71_n278_c;
                stage2_col72[6] = fa_s1_c71_n279_c;
                stage2_col72[7] = fa_s1_c72_n280_s;
                stage2_col72[8] = fa_s1_c72_n281_s;
                stage2_col72[9] = fa_s1_c72_n282_s;
                stage2_col72[10] = fa_s1_c72_n283_s;
                stage2_col72[11] = fa_s1_c72_n284_s;
                stage2_col72[12] = fa_s1_c72_n285_s;
                stage2_col72[13] = fa_s1_c72_n286_s;
                stage2_col73[0] = fa_s1_c72_n280_c;
                stage2_col73[1] = fa_s1_c72_n281_c;
                stage2_col73[2] = fa_s1_c72_n282_c;
                stage2_col73[3] = fa_s1_c72_n283_c;
                stage2_col73[4] = fa_s1_c72_n284_c;
                stage2_col73[5] = fa_s1_c72_n285_c;
                stage2_col73[6] = fa_s1_c72_n286_c;
                stage2_col73[7] = fa_s1_c73_n287_s;
                stage2_col73[8] = fa_s1_c73_n288_s;
                stage2_col73[9] = fa_s1_c73_n289_s;
                stage2_col73[10] = fa_s1_c73_n290_s;
                stage2_col73[11] = fa_s1_c73_n291_s;
                stage2_col73[12] = fa_s1_c73_n292_s;
                stage2_col73[13] = fa_s1_c73_n293_s;
                stage2_col73[14] = stage1_col73[21];
                stage2_col73[15] = stage1_col73[22];
                stage2_col74[0] = fa_s1_c73_n287_c;
                stage2_col74[1] = fa_s1_c73_n288_c;
                stage2_col74[2] = fa_s1_c73_n289_c;
                stage2_col74[3] = fa_s1_c73_n290_c;
                stage2_col74[4] = fa_s1_c73_n291_c;
                stage2_col74[5] = fa_s1_c73_n292_c;
                stage2_col74[6] = fa_s1_c73_n293_c;
                stage2_col74[7] = fa_s1_c74_n294_s;
                stage2_col74[8] = fa_s1_c74_n295_s;
                stage2_col74[9] = fa_s1_c74_n296_s;
                stage2_col74[10] = fa_s1_c74_n297_s;
                stage2_col74[11] = fa_s1_c74_n298_s;
                stage2_col74[12] = fa_s1_c74_n299_s;
                stage2_col74[13] = fa_s1_c74_n300_s;
                stage2_col75[0] = fa_s1_c74_n294_c;
                stage2_col75[1] = fa_s1_c74_n295_c;
                stage2_col75[2] = fa_s1_c74_n296_c;
                stage2_col75[3] = fa_s1_c74_n297_c;
                stage2_col75[4] = fa_s1_c74_n298_c;
                stage2_col75[5] = fa_s1_c74_n299_c;
                stage2_col75[6] = fa_s1_c74_n300_c;
                stage2_col75[7] = fa_s1_c75_n301_s;
                stage2_col75[8] = fa_s1_c75_n302_s;
                stage2_col75[9] = fa_s1_c75_n303_s;
                stage2_col75[10] = fa_s1_c75_n304_s;
                stage2_col75[11] = fa_s1_c75_n305_s;
                stage2_col75[12] = fa_s1_c75_n306_s;
                stage2_col75[13] = fa_s1_c75_n307_s;
                stage2_col75[14] = stage1_col75[21];
                stage2_col75[15] = stage1_col75[22];
                stage2_col76[0] = fa_s1_c75_n301_c;
                stage2_col76[1] = fa_s1_c75_n302_c;
                stage2_col76[2] = fa_s1_c75_n303_c;
                stage2_col76[3] = fa_s1_c75_n304_c;
                stage2_col76[4] = fa_s1_c75_n305_c;
                stage2_col76[5] = fa_s1_c75_n306_c;
                stage2_col76[6] = fa_s1_c75_n307_c;
                stage2_col76[7] = fa_s1_c76_n308_s;
                stage2_col76[8] = fa_s1_c76_n309_s;
                stage2_col76[9] = fa_s1_c76_n310_s;
                stage2_col76[10] = fa_s1_c76_n311_s;
                stage2_col76[11] = fa_s1_c76_n312_s;
                stage2_col76[12] = fa_s1_c76_n313_s;
                stage2_col76[13] = fa_s1_c76_n314_s;
                stage2_col77[0] = fa_s1_c76_n308_c;
                stage2_col77[1] = fa_s1_c76_n309_c;
                stage2_col77[2] = fa_s1_c76_n310_c;
                stage2_col77[3] = fa_s1_c76_n311_c;
                stage2_col77[4] = fa_s1_c76_n312_c;
                stage2_col77[5] = fa_s1_c76_n313_c;
                stage2_col77[6] = fa_s1_c76_n314_c;
                stage2_col77[7] = fa_s1_c77_n315_s;
                stage2_col77[8] = fa_s1_c77_n316_s;
                stage2_col77[9] = fa_s1_c77_n317_s;
                stage2_col77[10] = fa_s1_c77_n318_s;
                stage2_col77[11] = fa_s1_c77_n319_s;
                stage2_col77[12] = fa_s1_c77_n320_s;
                stage2_col77[13] = fa_s1_c77_n321_s;
                stage2_col77[14] = stage1_col77[21];
                stage2_col77[15] = stage1_col77[22];
                stage2_col78[0] = fa_s1_c77_n315_c;
                stage2_col78[1] = fa_s1_c77_n316_c;
                stage2_col78[2] = fa_s1_c77_n317_c;
                stage2_col78[3] = fa_s1_c77_n318_c;
                stage2_col78[4] = fa_s1_c77_n319_c;
                stage2_col78[5] = fa_s1_c77_n320_c;
                stage2_col78[6] = fa_s1_c77_n321_c;
                stage2_col78[7] = fa_s1_c78_n322_s;
                stage2_col78[8] = fa_s1_c78_n323_s;
                stage2_col78[9] = fa_s1_c78_n324_s;
                stage2_col78[10] = fa_s1_c78_n325_s;
                stage2_col78[11] = fa_s1_c78_n326_s;
                stage2_col78[12] = fa_s1_c78_n327_s;
                stage2_col78[13] = fa_s1_c78_n328_s;
                stage2_col79[0] = fa_s1_c78_n322_c;
                stage2_col79[1] = fa_s1_c78_n323_c;
                stage2_col79[2] = fa_s1_c78_n324_c;
                stage2_col79[3] = fa_s1_c78_n325_c;
                stage2_col79[4] = fa_s1_c78_n326_c;
                stage2_col79[5] = fa_s1_c78_n327_c;
                stage2_col79[6] = fa_s1_c78_n328_c;
                stage2_col79[7] = fa_s1_c79_n329_s;
                stage2_col79[8] = fa_s1_c79_n330_s;
                stage2_col79[9] = fa_s1_c79_n331_s;
                stage2_col79[10] = fa_s1_c79_n332_s;
                stage2_col79[11] = fa_s1_c79_n333_s;
                stage2_col79[12] = fa_s1_c79_n334_s;
                stage2_col79[13] = fa_s1_c79_n335_s;
                stage2_col79[14] = stage1_col79[21];
                stage2_col79[15] = stage1_col79[22];
                stage2_col80[0] = fa_s1_c79_n329_c;
                stage2_col80[1] = fa_s1_c79_n330_c;
                stage2_col80[2] = fa_s1_c79_n331_c;
                stage2_col80[3] = fa_s1_c79_n332_c;
                stage2_col80[4] = fa_s1_c79_n333_c;
                stage2_col80[5] = fa_s1_c79_n334_c;
                stage2_col80[6] = fa_s1_c79_n335_c;
                stage2_col80[7] = fa_s1_c80_n336_s;
                stage2_col80[8] = fa_s1_c80_n337_s;
                stage2_col80[9] = fa_s1_c80_n338_s;
                stage2_col80[10] = fa_s1_c80_n339_s;
                stage2_col80[11] = fa_s1_c80_n340_s;
                stage2_col80[12] = fa_s1_c80_n341_s;
                stage2_col80[13] = fa_s1_c80_n342_s;
                stage2_col81[0] = fa_s1_c80_n336_c;
                stage2_col81[1] = fa_s1_c80_n337_c;
                stage2_col81[2] = fa_s1_c80_n338_c;
                stage2_col81[3] = fa_s1_c80_n339_c;
                stage2_col81[4] = fa_s1_c80_n340_c;
                stage2_col81[5] = fa_s1_c80_n341_c;
                stage2_col81[6] = fa_s1_c80_n342_c;
                stage2_col81[7] = fa_s1_c81_n343_s;
                stage2_col81[8] = fa_s1_c81_n344_s;
                stage2_col81[9] = fa_s1_c81_n345_s;
                stage2_col81[10] = fa_s1_c81_n346_s;
                stage2_col81[11] = fa_s1_c81_n347_s;
                stage2_col81[12] = fa_s1_c81_n348_s;
                stage2_col81[13] = fa_s1_c81_n349_s;
                stage2_col81[14] = stage1_col81[21];
                stage2_col81[15] = stage1_col81[22];
                stage2_col82[0] = fa_s1_c81_n343_c;
                stage2_col82[1] = fa_s1_c81_n344_c;
                stage2_col82[2] = fa_s1_c81_n345_c;
                stage2_col82[3] = fa_s1_c81_n346_c;
                stage2_col82[4] = fa_s1_c81_n347_c;
                stage2_col82[5] = fa_s1_c81_n348_c;
                stage2_col82[6] = fa_s1_c81_n349_c;
                stage2_col82[7] = fa_s1_c82_n350_s;
                stage2_col82[8] = fa_s1_c82_n351_s;
                stage2_col82[9] = fa_s1_c82_n352_s;
                stage2_col82[10] = fa_s1_c82_n353_s;
                stage2_col82[11] = fa_s1_c82_n354_s;
                stage2_col82[12] = fa_s1_c82_n355_s;
                stage2_col82[13] = fa_s1_c82_n356_s;
                stage2_col83[0] = fa_s1_c82_n350_c;
                stage2_col83[1] = fa_s1_c82_n351_c;
                stage2_col83[2] = fa_s1_c82_n352_c;
                stage2_col83[3] = fa_s1_c82_n353_c;
                stage2_col83[4] = fa_s1_c82_n354_c;
                stage2_col83[5] = fa_s1_c82_n355_c;
                stage2_col83[6] = fa_s1_c82_n356_c;
                stage2_col83[7] = fa_s1_c83_n357_s;
                stage2_col83[8] = fa_s1_c83_n358_s;
                stage2_col83[9] = fa_s1_c83_n359_s;
                stage2_col83[10] = fa_s1_c83_n360_s;
                stage2_col83[11] = fa_s1_c83_n361_s;
                stage2_col83[12] = fa_s1_c83_n362_s;
                stage2_col83[13] = fa_s1_c83_n363_s;
                stage2_col83[14] = stage1_col83[21];
                stage2_col83[15] = stage1_col83[22];
                stage2_col84[0] = fa_s1_c83_n357_c;
                stage2_col84[1] = fa_s1_c83_n358_c;
                stage2_col84[2] = fa_s1_c83_n359_c;
                stage2_col84[3] = fa_s1_c83_n360_c;
                stage2_col84[4] = fa_s1_c83_n361_c;
                stage2_col84[5] = fa_s1_c83_n362_c;
                stage2_col84[6] = fa_s1_c83_n363_c;
                stage2_col84[7] = fa_s1_c84_n364_s;
                stage2_col84[8] = fa_s1_c84_n365_s;
                stage2_col84[9] = fa_s1_c84_n366_s;
                stage2_col84[10] = fa_s1_c84_n367_s;
                stage2_col84[11] = fa_s1_c84_n368_s;
                stage2_col84[12] = fa_s1_c84_n369_s;
                stage2_col84[13] = fa_s1_c84_n370_s;
                stage2_col85[0] = fa_s1_c84_n364_c;
                stage2_col85[1] = fa_s1_c84_n365_c;
                stage2_col85[2] = fa_s1_c84_n366_c;
                stage2_col85[3] = fa_s1_c84_n367_c;
                stage2_col85[4] = fa_s1_c84_n368_c;
                stage2_col85[5] = fa_s1_c84_n369_c;
                stage2_col85[6] = fa_s1_c84_n370_c;
                stage2_col85[7] = fa_s1_c85_n371_s;
                stage2_col85[8] = fa_s1_c85_n372_s;
                stage2_col85[9] = fa_s1_c85_n373_s;
                stage2_col85[10] = fa_s1_c85_n374_s;
                stage2_col85[11] = fa_s1_c85_n375_s;
                stage2_col85[12] = fa_s1_c85_n376_s;
                stage2_col85[13] = fa_s1_c85_n377_s;
                stage2_col85[14] = stage1_col85[21];
                stage2_col85[15] = stage1_col85[22];
                stage2_col86[0] = fa_s1_c85_n371_c;
                stage2_col86[1] = fa_s1_c85_n372_c;
                stage2_col86[2] = fa_s1_c85_n373_c;
                stage2_col86[3] = fa_s1_c85_n374_c;
                stage2_col86[4] = fa_s1_c85_n375_c;
                stage2_col86[5] = fa_s1_c85_n376_c;
                stage2_col86[6] = fa_s1_c85_n377_c;
                stage2_col86[7] = fa_s1_c86_n378_s;
                stage2_col86[8] = fa_s1_c86_n379_s;
                stage2_col86[9] = fa_s1_c86_n380_s;
                stage2_col86[10] = fa_s1_c86_n381_s;
                stage2_col86[11] = fa_s1_c86_n382_s;
                stage2_col86[12] = fa_s1_c86_n383_s;
                stage2_col86[13] = fa_s1_c86_n384_s;
                stage2_col87[0] = fa_s1_c86_n378_c;
                stage2_col87[1] = fa_s1_c86_n379_c;
                stage2_col87[2] = fa_s1_c86_n380_c;
                stage2_col87[3] = fa_s1_c86_n381_c;
                stage2_col87[4] = fa_s1_c86_n382_c;
                stage2_col87[5] = fa_s1_c86_n383_c;
                stage2_col87[6] = fa_s1_c86_n384_c;
                stage2_col87[7] = fa_s1_c87_n385_s;
                stage2_col87[8] = fa_s1_c87_n386_s;
                stage2_col87[9] = fa_s1_c87_n387_s;
                stage2_col87[10] = fa_s1_c87_n388_s;
                stage2_col87[11] = fa_s1_c87_n389_s;
                stage2_col87[12] = fa_s1_c87_n390_s;
                stage2_col87[13] = fa_s1_c87_n391_s;
                stage2_col87[14] = stage1_col87[21];
                stage2_col87[15] = stage1_col87[22];
                stage2_col88[0] = fa_s1_c87_n385_c;
                stage2_col88[1] = fa_s1_c87_n386_c;
                stage2_col88[2] = fa_s1_c87_n387_c;
                stage2_col88[3] = fa_s1_c87_n388_c;
                stage2_col88[4] = fa_s1_c87_n389_c;
                stage2_col88[5] = fa_s1_c87_n390_c;
                stage2_col88[6] = fa_s1_c87_n391_c;
                stage2_col88[7] = fa_s1_c88_n392_s;
                stage2_col88[8] = fa_s1_c88_n393_s;
                stage2_col88[9] = fa_s1_c88_n394_s;
                stage2_col88[10] = fa_s1_c88_n395_s;
                stage2_col88[11] = fa_s1_c88_n396_s;
                stage2_col88[12] = fa_s1_c88_n397_s;
                stage2_col88[13] = fa_s1_c88_n398_s;
                stage2_col89[0] = fa_s1_c88_n392_c;
                stage2_col89[1] = fa_s1_c88_n393_c;
                stage2_col89[2] = fa_s1_c88_n394_c;
                stage2_col89[3] = fa_s1_c88_n395_c;
                stage2_col89[4] = fa_s1_c88_n396_c;
                stage2_col89[5] = fa_s1_c88_n397_c;
                stage2_col89[6] = fa_s1_c88_n398_c;
                stage2_col89[7] = fa_s1_c89_n399_s;
                stage2_col89[8] = fa_s1_c89_n400_s;
                stage2_col89[9] = fa_s1_c89_n401_s;
                stage2_col89[10] = fa_s1_c89_n402_s;
                stage2_col89[11] = fa_s1_c89_n403_s;
                stage2_col89[12] = fa_s1_c89_n404_s;
                stage2_col89[13] = fa_s1_c89_n405_s;
                stage2_col89[14] = stage1_col89[21];
                stage2_col89[15] = stage1_col89[22];
                stage2_col90[0] = fa_s1_c89_n399_c;
                stage2_col90[1] = fa_s1_c89_n400_c;
                stage2_col90[2] = fa_s1_c89_n401_c;
                stage2_col90[3] = fa_s1_c89_n402_c;
                stage2_col90[4] = fa_s1_c89_n403_c;
                stage2_col90[5] = fa_s1_c89_n404_c;
                stage2_col90[6] = fa_s1_c89_n405_c;
                stage2_col90[7] = fa_s1_c90_n406_s;
                stage2_col90[8] = fa_s1_c90_n407_s;
                stage2_col90[9] = fa_s1_c90_n408_s;
                stage2_col90[10] = fa_s1_c90_n409_s;
                stage2_col90[11] = fa_s1_c90_n410_s;
                stage2_col90[12] = fa_s1_c90_n411_s;
                stage2_col90[13] = fa_s1_c90_n412_s;
                stage2_col91[0] = fa_s1_c90_n406_c;
                stage2_col91[1] = fa_s1_c90_n407_c;
                stage2_col91[2] = fa_s1_c90_n408_c;
                stage2_col91[3] = fa_s1_c90_n409_c;
                stage2_col91[4] = fa_s1_c90_n410_c;
                stage2_col91[5] = fa_s1_c90_n411_c;
                stage2_col91[6] = fa_s1_c90_n412_c;
                stage2_col91[7] = fa_s1_c91_n413_s;
                stage2_col91[8] = fa_s1_c91_n414_s;
                stage2_col91[9] = fa_s1_c91_n415_s;
                stage2_col91[10] = fa_s1_c91_n416_s;
                stage2_col91[11] = fa_s1_c91_n417_s;
                stage2_col91[12] = fa_s1_c91_n418_s;
                stage2_col91[13] = fa_s1_c91_n419_s;
                stage2_col91[14] = stage1_col91[21];
                stage2_col91[15] = stage1_col91[22];
                stage2_col92[0] = fa_s1_c91_n413_c;
                stage2_col92[1] = fa_s1_c91_n414_c;
                stage2_col92[2] = fa_s1_c91_n415_c;
                stage2_col92[3] = fa_s1_c91_n416_c;
                stage2_col92[4] = fa_s1_c91_n417_c;
                stage2_col92[5] = fa_s1_c91_n418_c;
                stage2_col92[6] = fa_s1_c91_n419_c;
                stage2_col92[7] = fa_s1_c92_n420_s;
                stage2_col92[8] = fa_s1_c92_n421_s;
                stage2_col92[9] = fa_s1_c92_n422_s;
                stage2_col92[10] = fa_s1_c92_n423_s;
                stage2_col92[11] = fa_s1_c92_n424_s;
                stage2_col92[12] = fa_s1_c92_n425_s;
                stage2_col92[13] = fa_s1_c92_n426_s;
                stage2_col93[0] = fa_s1_c92_n420_c;
                stage2_col93[1] = fa_s1_c92_n421_c;
                stage2_col93[2] = fa_s1_c92_n422_c;
                stage2_col93[3] = fa_s1_c92_n423_c;
                stage2_col93[4] = fa_s1_c92_n424_c;
                stage2_col93[5] = fa_s1_c92_n425_c;
                stage2_col93[6] = fa_s1_c92_n426_c;
                stage2_col93[7] = fa_s1_c93_n427_s;
                stage2_col93[8] = fa_s1_c93_n428_s;
                stage2_col93[9] = fa_s1_c93_n429_s;
                stage2_col93[10] = fa_s1_c93_n430_s;
                stage2_col93[11] = fa_s1_c93_n431_s;
                stage2_col93[12] = fa_s1_c93_n432_s;
                stage2_col93[13] = fa_s1_c93_n433_s;
                stage2_col93[14] = stage1_col93[21];
                stage2_col93[15] = stage1_col93[22];
                stage2_col94[0] = fa_s1_c93_n427_c;
                stage2_col94[1] = fa_s1_c93_n428_c;
                stage2_col94[2] = fa_s1_c93_n429_c;
                stage2_col94[3] = fa_s1_c93_n430_c;
                stage2_col94[4] = fa_s1_c93_n431_c;
                stage2_col94[5] = fa_s1_c93_n432_c;
                stage2_col94[6] = fa_s1_c93_n433_c;
                stage2_col94[7] = fa_s1_c94_n434_s;
                stage2_col94[8] = fa_s1_c94_n435_s;
                stage2_col94[9] = fa_s1_c94_n436_s;
                stage2_col94[10] = fa_s1_c94_n437_s;
                stage2_col94[11] = fa_s1_c94_n438_s;
                stage2_col94[12] = fa_s1_c94_n439_s;
                stage2_col94[13] = fa_s1_c94_n440_s;
                stage2_col95[0] = fa_s1_c94_n434_c;
                stage2_col95[1] = fa_s1_c94_n435_c;
                stage2_col95[2] = fa_s1_c94_n436_c;
                stage2_col95[3] = fa_s1_c94_n437_c;
                stage2_col95[4] = fa_s1_c94_n438_c;
                stage2_col95[5] = fa_s1_c94_n439_c;
                stage2_col95[6] = fa_s1_c94_n440_c;
                stage2_col95[7] = fa_s1_c95_n441_s;
                stage2_col95[8] = fa_s1_c95_n442_s;
                stage2_col95[9] = fa_s1_c95_n443_s;
                stage2_col95[10] = fa_s1_c95_n444_s;
                stage2_col95[11] = fa_s1_c95_n445_s;
                stage2_col95[12] = fa_s1_c95_n446_s;
                stage2_col95[13] = fa_s1_c95_n447_s;
                stage2_col95[14] = stage1_col95[21];
                stage2_col95[15] = stage1_col95[22];
                stage2_col96[0] = fa_s1_c95_n441_c;
                stage2_col96[1] = fa_s1_c95_n442_c;
                stage2_col96[2] = fa_s1_c95_n443_c;
                stage2_col96[3] = fa_s1_c95_n444_c;
                stage2_col96[4] = fa_s1_c95_n445_c;
                stage2_col96[5] = fa_s1_c95_n446_c;
                stage2_col96[6] = fa_s1_c95_n447_c;
                stage2_col96[7] = fa_s1_c96_n448_s;
                stage2_col96[8] = fa_s1_c96_n449_s;
                stage2_col96[9] = fa_s1_c96_n450_s;
                stage2_col96[10] = fa_s1_c96_n451_s;
                stage2_col96[11] = fa_s1_c96_n452_s;
                stage2_col96[12] = fa_s1_c96_n453_s;
                stage2_col96[13] = fa_s1_c96_n454_s;
                stage2_col97[0] = fa_s1_c96_n448_c;
                stage2_col97[1] = fa_s1_c96_n449_c;
                stage2_col97[2] = fa_s1_c96_n450_c;
                stage2_col97[3] = fa_s1_c96_n451_c;
                stage2_col97[4] = fa_s1_c96_n452_c;
                stage2_col97[5] = fa_s1_c96_n453_c;
                stage2_col97[6] = fa_s1_c96_n454_c;
                stage2_col97[7] = fa_s1_c97_n455_s;
                stage2_col97[8] = fa_s1_c97_n456_s;
                stage2_col97[9] = fa_s1_c97_n457_s;
                stage2_col97[10] = fa_s1_c97_n458_s;
                stage2_col97[11] = fa_s1_c97_n459_s;
                stage2_col97[12] = fa_s1_c97_n460_s;
                stage2_col97[13] = fa_s1_c97_n461_s;
                stage2_col97[14] = stage1_col97[21];
                stage2_col97[15] = stage1_col97[22];
                stage2_col98[0] = fa_s1_c97_n455_c;
                stage2_col98[1] = fa_s1_c97_n456_c;
                stage2_col98[2] = fa_s1_c97_n457_c;
                stage2_col98[3] = fa_s1_c97_n458_c;
                stage2_col98[4] = fa_s1_c97_n459_c;
                stage2_col98[5] = fa_s1_c97_n460_c;
                stage2_col98[6] = fa_s1_c97_n461_c;
                stage2_col98[7] = fa_s1_c98_n462_s;
                stage2_col98[8] = fa_s1_c98_n463_s;
                stage2_col98[9] = fa_s1_c98_n464_s;
                stage2_col98[10] = fa_s1_c98_n465_s;
                stage2_col98[11] = fa_s1_c98_n466_s;
                stage2_col98[12] = fa_s1_c98_n467_s;
                stage2_col98[13] = fa_s1_c98_n468_s;
                stage2_col99[0] = fa_s1_c98_n462_c;
                stage2_col99[1] = fa_s1_c98_n463_c;
                stage2_col99[2] = fa_s1_c98_n464_c;
                stage2_col99[3] = fa_s1_c98_n465_c;
                stage2_col99[4] = fa_s1_c98_n466_c;
                stage2_col99[5] = fa_s1_c98_n467_c;
                stage2_col99[6] = fa_s1_c98_n468_c;
                stage2_col99[7] = fa_s1_c99_n469_s;
                stage2_col99[8] = fa_s1_c99_n470_s;
                stage2_col99[9] = fa_s1_c99_n471_s;
                stage2_col99[10] = fa_s1_c99_n472_s;
                stage2_col99[11] = fa_s1_c99_n473_s;
                stage2_col99[12] = fa_s1_c99_n474_s;
                stage2_col99[13] = fa_s1_c99_n475_s;
                stage2_col99[14] = stage1_col99[21];
                stage2_col99[15] = stage1_col99[22];
                stage2_col100[0] = fa_s1_c99_n469_c;
                stage2_col100[1] = fa_s1_c99_n470_c;
                stage2_col100[2] = fa_s1_c99_n471_c;
                stage2_col100[3] = fa_s1_c99_n472_c;
                stage2_col100[4] = fa_s1_c99_n473_c;
                stage2_col100[5] = fa_s1_c99_n474_c;
                stage2_col100[6] = fa_s1_c99_n475_c;
                stage2_col100[7] = fa_s1_c100_n476_s;
                stage2_col100[8] = fa_s1_c100_n477_s;
                stage2_col100[9] = fa_s1_c100_n478_s;
                stage2_col100[10] = fa_s1_c100_n479_s;
                stage2_col100[11] = fa_s1_c100_n480_s;
                stage2_col100[12] = fa_s1_c100_n481_s;
                stage2_col100[13] = fa_s1_c100_n482_s;
                stage2_col101[0] = fa_s1_c100_n476_c;
                stage2_col101[1] = fa_s1_c100_n477_c;
                stage2_col101[2] = fa_s1_c100_n478_c;
                stage2_col101[3] = fa_s1_c100_n479_c;
                stage2_col101[4] = fa_s1_c100_n480_c;
                stage2_col101[5] = fa_s1_c100_n481_c;
                stage2_col101[6] = fa_s1_c100_n482_c;
                stage2_col101[7] = fa_s1_c101_n483_s;
                stage2_col101[8] = fa_s1_c101_n484_s;
                stage2_col101[9] = fa_s1_c101_n485_s;
                stage2_col101[10] = fa_s1_c101_n486_s;
                stage2_col101[11] = fa_s1_c101_n487_s;
                stage2_col101[12] = fa_s1_c101_n488_s;
                stage2_col101[13] = fa_s1_c101_n489_s;
                stage2_col101[14] = stage1_col101[21];
                stage2_col101[15] = stage1_col101[22];
                stage2_col102[0] = fa_s1_c101_n483_c;
                stage2_col102[1] = fa_s1_c101_n484_c;
                stage2_col102[2] = fa_s1_c101_n485_c;
                stage2_col102[3] = fa_s1_c101_n486_c;
                stage2_col102[4] = fa_s1_c101_n487_c;
                stage2_col102[5] = fa_s1_c101_n488_c;
                stage2_col102[6] = fa_s1_c101_n489_c;
                stage2_col102[7] = fa_s1_c102_n490_s;
                stage2_col102[8] = fa_s1_c102_n491_s;
                stage2_col102[9] = fa_s1_c102_n492_s;
                stage2_col102[10] = fa_s1_c102_n493_s;
                stage2_col102[11] = fa_s1_c102_n494_s;
                stage2_col102[12] = fa_s1_c102_n495_s;
                stage2_col102[13] = fa_s1_c102_n496_s;
                stage2_col103[0] = fa_s1_c102_n490_c;
                stage2_col103[1] = fa_s1_c102_n491_c;
                stage2_col103[2] = fa_s1_c102_n492_c;
                stage2_col103[3] = fa_s1_c102_n493_c;
                stage2_col103[4] = fa_s1_c102_n494_c;
                stage2_col103[5] = fa_s1_c102_n495_c;
                stage2_col103[6] = fa_s1_c102_n496_c;
                stage2_col103[7] = fa_s1_c103_n497_s;
                stage2_col103[8] = fa_s1_c103_n498_s;
                stage2_col103[9] = fa_s1_c103_n499_s;
                stage2_col103[10] = fa_s1_c103_n500_s;
                stage2_col103[11] = fa_s1_c103_n501_s;
                stage2_col103[12] = fa_s1_c103_n502_s;
                stage2_col103[13] = fa_s1_c103_n503_s;
                stage2_col103[14] = stage1_col103[21];
                stage2_col103[15] = stage1_col103[22];
                stage2_col104[0] = fa_s1_c103_n497_c;
                stage2_col104[1] = fa_s1_c103_n498_c;
                stage2_col104[2] = fa_s1_c103_n499_c;
                stage2_col104[3] = fa_s1_c103_n500_c;
                stage2_col104[4] = fa_s1_c103_n501_c;
                stage2_col104[5] = fa_s1_c103_n502_c;
                stage2_col104[6] = fa_s1_c103_n503_c;
                stage2_col104[7] = fa_s1_c104_n504_s;
                stage2_col104[8] = fa_s1_c104_n505_s;
                stage2_col104[9] = fa_s1_c104_n506_s;
                stage2_col104[10] = fa_s1_c104_n507_s;
                stage2_col104[11] = fa_s1_c104_n508_s;
                stage2_col104[12] = fa_s1_c104_n509_s;
                stage2_col104[13] = fa_s1_c104_n510_s;
                stage2_col105[0] = fa_s1_c104_n504_c;
                stage2_col105[1] = fa_s1_c104_n505_c;
                stage2_col105[2] = fa_s1_c104_n506_c;
                stage2_col105[3] = fa_s1_c104_n507_c;
                stage2_col105[4] = fa_s1_c104_n508_c;
                stage2_col105[5] = fa_s1_c104_n509_c;
                stage2_col105[6] = fa_s1_c104_n510_c;
                stage2_col105[7] = fa_s1_c105_n511_s;
                stage2_col105[8] = fa_s1_c105_n512_s;
                stage2_col105[9] = fa_s1_c105_n513_s;
                stage2_col105[10] = fa_s1_c105_n514_s;
                stage2_col105[11] = fa_s1_c105_n515_s;
                stage2_col105[12] = fa_s1_c105_n516_s;
                stage2_col105[13] = fa_s1_c105_n517_s;
                stage2_col105[14] = stage1_col105[21];
                stage2_col105[15] = stage1_col105[22];
                stage2_col106[0] = fa_s1_c105_n511_c;
                stage2_col106[1] = fa_s1_c105_n512_c;
                stage2_col106[2] = fa_s1_c105_n513_c;
                stage2_col106[3] = fa_s1_c105_n514_c;
                stage2_col106[4] = fa_s1_c105_n515_c;
                stage2_col106[5] = fa_s1_c105_n516_c;
                stage2_col106[6] = fa_s1_c105_n517_c;
                stage2_col106[7] = fa_s1_c106_n518_s;
                stage2_col106[8] = fa_s1_c106_n519_s;
                stage2_col106[9] = fa_s1_c106_n520_s;
                stage2_col106[10] = fa_s1_c106_n521_s;
                stage2_col106[11] = fa_s1_c106_n522_s;
                stage2_col106[12] = fa_s1_c106_n523_s;
                stage2_col106[13] = fa_s1_c106_n524_s;
                stage2_col107[0] = fa_s1_c106_n518_c;
                stage2_col107[1] = fa_s1_c106_n519_c;
                stage2_col107[2] = fa_s1_c106_n520_c;
                stage2_col107[3] = fa_s1_c106_n521_c;
                stage2_col107[4] = fa_s1_c106_n522_c;
                stage2_col107[5] = fa_s1_c106_n523_c;
                stage2_col107[6] = fa_s1_c106_n524_c;
                stage2_col107[7] = fa_s1_c107_n525_s;
                stage2_col107[8] = fa_s1_c107_n526_s;
                stage2_col107[9] = fa_s1_c107_n527_s;
                stage2_col107[10] = fa_s1_c107_n528_s;
                stage2_col107[11] = fa_s1_c107_n529_s;
                stage2_col107[12] = fa_s1_c107_n530_s;
                stage2_col107[13] = fa_s1_c107_n531_s;
                stage2_col107[14] = stage1_col107[21];
                stage2_col107[15] = stage1_col107[22];
                stage2_col108[0] = fa_s1_c107_n525_c;
                stage2_col108[1] = fa_s1_c107_n526_c;
                stage2_col108[2] = fa_s1_c107_n527_c;
                stage2_col108[3] = fa_s1_c107_n528_c;
                stage2_col108[4] = fa_s1_c107_n529_c;
                stage2_col108[5] = fa_s1_c107_n530_c;
                stage2_col108[6] = fa_s1_c107_n531_c;
                stage2_col108[7] = fa_s1_c108_n532_s;
                stage2_col108[8] = fa_s1_c108_n533_s;
                stage2_col108[9] = fa_s1_c108_n534_s;
                stage2_col108[10] = fa_s1_c108_n535_s;
                stage2_col108[11] = fa_s1_c108_n536_s;
                stage2_col108[12] = fa_s1_c108_n537_s;
                stage2_col108[13] = fa_s1_c108_n538_s;
                stage2_col109[0] = fa_s1_c108_n532_c;
                stage2_col109[1] = fa_s1_c108_n533_c;
                stage2_col109[2] = fa_s1_c108_n534_c;
                stage2_col109[3] = fa_s1_c108_n535_c;
                stage2_col109[4] = fa_s1_c108_n536_c;
                stage2_col109[5] = fa_s1_c108_n537_c;
                stage2_col109[6] = fa_s1_c108_n538_c;
                stage2_col109[7] = fa_s1_c109_n539_s;
                stage2_col109[8] = fa_s1_c109_n540_s;
                stage2_col109[9] = fa_s1_c109_n541_s;
                stage2_col109[10] = fa_s1_c109_n542_s;
                stage2_col109[11] = fa_s1_c109_n543_s;
                stage2_col109[12] = fa_s1_c109_n544_s;
                stage2_col109[13] = fa_s1_c109_n545_s;
                stage2_col109[14] = stage1_col109[21];
                stage2_col109[15] = stage1_col109[22];
                stage2_col110[0] = fa_s1_c109_n539_c;
                stage2_col110[1] = fa_s1_c109_n540_c;
                stage2_col110[2] = fa_s1_c109_n541_c;
                stage2_col110[3] = fa_s1_c109_n542_c;
                stage2_col110[4] = fa_s1_c109_n543_c;
                stage2_col110[5] = fa_s1_c109_n544_c;
                stage2_col110[6] = fa_s1_c109_n545_c;
                stage2_col110[7] = fa_s1_c110_n546_s;
                stage2_col110[8] = fa_s1_c110_n547_s;
                stage2_col110[9] = fa_s1_c110_n548_s;
                stage2_col110[10] = fa_s1_c110_n549_s;
                stage2_col110[11] = fa_s1_c110_n550_s;
                stage2_col110[12] = fa_s1_c110_n551_s;
                stage2_col110[13] = fa_s1_c110_n552_s;
                stage2_col111[0] = fa_s1_c110_n546_c;
                stage2_col111[1] = fa_s1_c110_n547_c;
                stage2_col111[2] = fa_s1_c110_n548_c;
                stage2_col111[3] = fa_s1_c110_n549_c;
                stage2_col111[4] = fa_s1_c110_n550_c;
                stage2_col111[5] = fa_s1_c110_n551_c;
                stage2_col111[6] = fa_s1_c110_n552_c;
                stage2_col111[7] = fa_s1_c111_n553_s;
                stage2_col111[8] = fa_s1_c111_n554_s;
                stage2_col111[9] = fa_s1_c111_n555_s;
                stage2_col111[10] = fa_s1_c111_n556_s;
                stage2_col111[11] = fa_s1_c111_n557_s;
                stage2_col111[12] = fa_s1_c111_n558_s;
                stage2_col111[13] = fa_s1_c111_n559_s;
                stage2_col111[14] = stage1_col111[21];
                stage2_col111[15] = stage1_col111[22];
                stage2_col112[0] = fa_s1_c111_n553_c;
                stage2_col112[1] = fa_s1_c111_n554_c;
                stage2_col112[2] = fa_s1_c111_n555_c;
                stage2_col112[3] = fa_s1_c111_n556_c;
                stage2_col112[4] = fa_s1_c111_n557_c;
                stage2_col112[5] = fa_s1_c111_n558_c;
                stage2_col112[6] = fa_s1_c111_n559_c;
                stage2_col112[7] = fa_s1_c112_n560_s;
                stage2_col112[8] = fa_s1_c112_n561_s;
                stage2_col112[9] = fa_s1_c112_n562_s;
                stage2_col112[10] = fa_s1_c112_n563_s;
                stage2_col112[11] = fa_s1_c112_n564_s;
                stage2_col112[12] = fa_s1_c112_n565_s;
                stage2_col112[13] = fa_s1_c112_n566_s;
                stage2_col113[0] = fa_s1_c112_n560_c;
                stage2_col113[1] = fa_s1_c112_n561_c;
                stage2_col113[2] = fa_s1_c112_n562_c;
                stage2_col113[3] = fa_s1_c112_n563_c;
                stage2_col113[4] = fa_s1_c112_n564_c;
                stage2_col113[5] = fa_s1_c112_n565_c;
                stage2_col113[6] = fa_s1_c112_n566_c;
                stage2_col113[7] = fa_s1_c113_n567_s;
                stage2_col113[8] = fa_s1_c113_n568_s;
                stage2_col113[9] = fa_s1_c113_n569_s;
                stage2_col113[10] = fa_s1_c113_n570_s;
                stage2_col113[11] = fa_s1_c113_n571_s;
                stage2_col113[12] = fa_s1_c113_n572_s;
                stage2_col113[13] = fa_s1_c113_n573_s;
                stage2_col113[14] = stage1_col113[21];
                stage2_col113[15] = stage1_col113[22];
                stage2_col114[0] = fa_s1_c113_n567_c;
                stage2_col114[1] = fa_s1_c113_n568_c;
                stage2_col114[2] = fa_s1_c113_n569_c;
                stage2_col114[3] = fa_s1_c113_n570_c;
                stage2_col114[4] = fa_s1_c113_n571_c;
                stage2_col114[5] = fa_s1_c113_n572_c;
                stage2_col114[6] = fa_s1_c113_n573_c;
                stage2_col114[7] = fa_s1_c114_n574_s;
                stage2_col114[8] = fa_s1_c114_n575_s;
                stage2_col114[9] = fa_s1_c114_n576_s;
                stage2_col114[10] = fa_s1_c114_n577_s;
                stage2_col114[11] = fa_s1_c114_n578_s;
                stage2_col114[12] = fa_s1_c114_n579_s;
                stage2_col114[13] = fa_s1_c114_n580_s;
                stage2_col115[0] = fa_s1_c114_n574_c;
                stage2_col115[1] = fa_s1_c114_n575_c;
                stage2_col115[2] = fa_s1_c114_n576_c;
                stage2_col115[3] = fa_s1_c114_n577_c;
                stage2_col115[4] = fa_s1_c114_n578_c;
                stage2_col115[5] = fa_s1_c114_n579_c;
                stage2_col115[6] = fa_s1_c114_n580_c;
                stage2_col115[7] = fa_s1_c115_n581_s;
                stage2_col115[8] = fa_s1_c115_n582_s;
                stage2_col115[9] = fa_s1_c115_n583_s;
                stage2_col115[10] = fa_s1_c115_n584_s;
                stage2_col115[11] = fa_s1_c115_n585_s;
                stage2_col115[12] = fa_s1_c115_n586_s;
                stage2_col115[13] = fa_s1_c115_n587_s;
                stage2_col115[14] = stage1_col115[21];
                stage2_col115[15] = stage1_col115[22];
                stage2_col116[0] = fa_s1_c115_n581_c;
                stage2_col116[1] = fa_s1_c115_n582_c;
                stage2_col116[2] = fa_s1_c115_n583_c;
                stage2_col116[3] = fa_s1_c115_n584_c;
                stage2_col116[4] = fa_s1_c115_n585_c;
                stage2_col116[5] = fa_s1_c115_n586_c;
                stage2_col116[6] = fa_s1_c115_n587_c;
                stage2_col116[7] = fa_s1_c116_n588_s;
                stage2_col116[8] = fa_s1_c116_n589_s;
                stage2_col116[9] = fa_s1_c116_n590_s;
                stage2_col116[10] = fa_s1_c116_n591_s;
                stage2_col116[11] = fa_s1_c116_n592_s;
                stage2_col116[12] = fa_s1_c116_n593_s;
                stage2_col116[13] = fa_s1_c116_n594_s;
                stage2_col117[0] = fa_s1_c116_n588_c;
                stage2_col117[1] = fa_s1_c116_n589_c;
                stage2_col117[2] = fa_s1_c116_n590_c;
                stage2_col117[3] = fa_s1_c116_n591_c;
                stage2_col117[4] = fa_s1_c116_n592_c;
                stage2_col117[5] = fa_s1_c116_n593_c;
                stage2_col117[6] = fa_s1_c116_n594_c;
                stage2_col117[7] = fa_s1_c117_n595_s;
                stage2_col117[8] = fa_s1_c117_n596_s;
                stage2_col117[9] = fa_s1_c117_n597_s;
                stage2_col117[10] = fa_s1_c117_n598_s;
                stage2_col117[11] = fa_s1_c117_n599_s;
                stage2_col117[12] = fa_s1_c117_n600_s;
                stage2_col117[13] = fa_s1_c117_n601_s;
                stage2_col117[14] = stage1_col117[21];
                stage2_col117[15] = stage1_col117[22];
                stage2_col118[0] = fa_s1_c117_n595_c;
                stage2_col118[1] = fa_s1_c117_n596_c;
                stage2_col118[2] = fa_s1_c117_n597_c;
                stage2_col118[3] = fa_s1_c117_n598_c;
                stage2_col118[4] = fa_s1_c117_n599_c;
                stage2_col118[5] = fa_s1_c117_n600_c;
                stage2_col118[6] = fa_s1_c117_n601_c;
                stage2_col118[7] = fa_s1_c118_n602_s;
                stage2_col118[8] = fa_s1_c118_n603_s;
                stage2_col118[9] = fa_s1_c118_n604_s;
                stage2_col118[10] = fa_s1_c118_n605_s;
                stage2_col118[11] = fa_s1_c118_n606_s;
                stage2_col118[12] = fa_s1_c118_n607_s;
                stage2_col118[13] = fa_s1_c118_n608_s;
                stage2_col119[0] = fa_s1_c118_n602_c;
                stage2_col119[1] = fa_s1_c118_n603_c;
                stage2_col119[2] = fa_s1_c118_n604_c;
                stage2_col119[3] = fa_s1_c118_n605_c;
                stage2_col119[4] = fa_s1_c118_n606_c;
                stage2_col119[5] = fa_s1_c118_n607_c;
                stage2_col119[6] = fa_s1_c118_n608_c;
                stage2_col119[7] = fa_s1_c119_n609_s;
                stage2_col119[8] = fa_s1_c119_n610_s;
                stage2_col119[9] = fa_s1_c119_n611_s;
                stage2_col119[10] = fa_s1_c119_n612_s;
                stage2_col119[11] = fa_s1_c119_n613_s;
                stage2_col119[12] = fa_s1_c119_n614_s;
                stage2_col119[13] = fa_s1_c119_n615_s;
                stage2_col119[14] = stage1_col119[21];
                stage2_col119[15] = stage1_col119[22];
                stage2_col120[0] = fa_s1_c119_n609_c;
                stage2_col120[1] = fa_s1_c119_n610_c;
                stage2_col120[2] = fa_s1_c119_n611_c;
                stage2_col120[3] = fa_s1_c119_n612_c;
                stage2_col120[4] = fa_s1_c119_n613_c;
                stage2_col120[5] = fa_s1_c119_n614_c;
                stage2_col120[6] = fa_s1_c119_n615_c;
                stage2_col120[7] = fa_s1_c120_n616_s;
                stage2_col120[8] = fa_s1_c120_n617_s;
                stage2_col120[9] = fa_s1_c120_n618_s;
                stage2_col120[10] = fa_s1_c120_n619_s;
                stage2_col120[11] = fa_s1_c120_n620_s;
                stage2_col120[12] = fa_s1_c120_n621_s;
                stage2_col120[13] = fa_s1_c120_n622_s;
                stage2_col121[0] = fa_s1_c120_n616_c;
                stage2_col121[1] = fa_s1_c120_n617_c;
                stage2_col121[2] = fa_s1_c120_n618_c;
                stage2_col121[3] = fa_s1_c120_n619_c;
                stage2_col121[4] = fa_s1_c120_n620_c;
                stage2_col121[5] = fa_s1_c120_n621_c;
                stage2_col121[6] = fa_s1_c120_n622_c;
                stage2_col121[7] = fa_s1_c121_n623_s;
                stage2_col121[8] = fa_s1_c121_n624_s;
                stage2_col121[9] = fa_s1_c121_n625_s;
                stage2_col121[10] = fa_s1_c121_n626_s;
                stage2_col121[11] = fa_s1_c121_n627_s;
                stage2_col121[12] = fa_s1_c121_n628_s;
                stage2_col121[13] = fa_s1_c121_n629_s;
                stage2_col121[14] = stage1_col121[21];
                stage2_col121[15] = stage1_col121[22];
                stage2_col122[0] = fa_s1_c121_n623_c;
                stage2_col122[1] = fa_s1_c121_n624_c;
                stage2_col122[2] = fa_s1_c121_n625_c;
                stage2_col122[3] = fa_s1_c121_n626_c;
                stage2_col122[4] = fa_s1_c121_n627_c;
                stage2_col122[5] = fa_s1_c121_n628_c;
                stage2_col122[6] = fa_s1_c121_n629_c;
                stage2_col122[7] = fa_s1_c122_n630_s;
                stage2_col122[8] = fa_s1_c122_n631_s;
                stage2_col122[9] = fa_s1_c122_n632_s;
                stage2_col122[10] = fa_s1_c122_n633_s;
                stage2_col122[11] = fa_s1_c122_n634_s;
                stage2_col122[12] = fa_s1_c122_n635_s;
                stage2_col122[13] = fa_s1_c122_n636_s;
                stage2_col123[0] = fa_s1_c122_n630_c;
                stage2_col123[1] = fa_s1_c122_n631_c;
                stage2_col123[2] = fa_s1_c122_n632_c;
                stage2_col123[3] = fa_s1_c122_n633_c;
                stage2_col123[4] = fa_s1_c122_n634_c;
                stage2_col123[5] = fa_s1_c122_n635_c;
                stage2_col123[6] = fa_s1_c122_n636_c;
                stage2_col123[7] = fa_s1_c123_n637_s;
                stage2_col123[8] = fa_s1_c123_n638_s;
                stage2_col123[9] = fa_s1_c123_n639_s;
                stage2_col123[10] = fa_s1_c123_n640_s;
                stage2_col123[11] = fa_s1_c123_n641_s;
                stage2_col123[12] = fa_s1_c123_n642_s;
                stage2_col123[13] = fa_s1_c123_n643_s;
                stage2_col123[14] = stage1_col123[21];
                stage2_col123[15] = stage1_col123[22];
                stage2_col124[0] = fa_s1_c123_n637_c;
                stage2_col124[1] = fa_s1_c123_n638_c;
                stage2_col124[2] = fa_s1_c123_n639_c;
                stage2_col124[3] = fa_s1_c123_n640_c;
                stage2_col124[4] = fa_s1_c123_n641_c;
                stage2_col124[5] = fa_s1_c123_n642_c;
                stage2_col124[6] = fa_s1_c123_n643_c;
                stage2_col124[7] = fa_s1_c124_n644_s;
                stage2_col124[8] = fa_s1_c124_n645_s;
                stage2_col124[9] = fa_s1_c124_n646_s;
                stage2_col124[10] = fa_s1_c124_n647_s;
                stage2_col124[11] = fa_s1_c124_n648_s;
                stage2_col124[12] = fa_s1_c124_n649_s;
                stage2_col124[13] = fa_s1_c124_n650_s;
                stage2_col125[0] = fa_s1_c124_n644_c;
                stage2_col125[1] = fa_s1_c124_n645_c;
                stage2_col125[2] = fa_s1_c124_n646_c;
                stage2_col125[3] = fa_s1_c124_n647_c;
                stage2_col125[4] = fa_s1_c124_n648_c;
                stage2_col125[5] = fa_s1_c124_n649_c;
                stage2_col125[6] = fa_s1_c124_n650_c;
                stage2_col125[7] = fa_s1_c125_n651_s;
                stage2_col125[8] = fa_s1_c125_n652_s;
                stage2_col125[9] = fa_s1_c125_n653_s;
                stage2_col125[10] = fa_s1_c125_n654_s;
                stage2_col125[11] = fa_s1_c125_n655_s;
                stage2_col125[12] = fa_s1_c125_n656_s;
                stage2_col125[13] = fa_s1_c125_n657_s;
                stage2_col125[14] = stage1_col125[21];
                stage2_col125[15] = stage1_col125[22];
                stage2_col126[0] = fa_s1_c125_n651_c;
                stage2_col126[1] = fa_s1_c125_n652_c;
                stage2_col126[2] = fa_s1_c125_n653_c;
                stage2_col126[3] = fa_s1_c125_n654_c;
                stage2_col126[4] = fa_s1_c125_n655_c;
                stage2_col126[5] = fa_s1_c125_n656_c;
                stage2_col126[6] = fa_s1_c125_n657_c;
                stage2_col126[7] = fa_s1_c126_n658_s;
                stage2_col126[8] = fa_s1_c126_n659_s;
                stage2_col126[9] = fa_s1_c126_n660_s;
                stage2_col126[10] = fa_s1_c126_n661_s;
                stage2_col126[11] = fa_s1_c126_n662_s;
                stage2_col126[12] = fa_s1_c126_n663_s;
                stage2_col126[13] = fa_s1_c126_n664_s;
                stage2_col127[0] = fa_s1_c126_n658_c;
                stage2_col127[1] = fa_s1_c126_n659_c;
                stage2_col127[2] = fa_s1_c126_n660_c;
                stage2_col127[3] = fa_s1_c126_n661_c;
                stage2_col127[4] = fa_s1_c126_n662_c;
                stage2_col127[5] = fa_s1_c126_n663_c;
                stage2_col127[6] = fa_s1_c126_n664_c;
                stage2_col127[7] = stage1_col127[0];
                stage2_col127[8] = stage1_col127[1];
                stage2_col127[9] = stage1_col127[2];
                stage2_col127[10] = stage1_col127[3];
                stage2_col127[11] = stage1_col127[4];
                stage2_col127[12] = stage1_col127[5];
                stage2_col127[13] = stage1_col127[6];
                stage2_col127[14] = stage1_col127[7];
                stage2_col127[15] = stage1_col127[8];
                stage2_col127[16] = stage1_col127[9];
                stage2_col127[17] = stage1_col127[10];
                stage2_col127[18] = stage1_col127[11];
                stage2_col127[19] = stage1_col127[11];
                stage2_col127[20] = stage1_col127[11];
                stage2_col127[21] = stage1_col127[11];
                stage2_col127[22] = stage1_col127[11];
                stage2_col127[23] = stage1_col127[11];
                stage2_col127[24] = stage1_col127[11];
                stage2_col127[25] = stage1_col127[11];
                stage2_col127[26] = stage1_col127[11];
                stage2_col127[27] = stage1_col127[11];
                stage2_col127[28] = stage1_col127[11];
                stage2_col127[29] = stage1_col127[11];
                stage2_col127[30] = stage1_col127[11];
                stage2_col127[31] = stage1_col127[11];
                stage2_col127[32] = stage1_col127[11];
                stage2_col127[33] = stage1_col127[11];
                stage2_col127[34] = stage1_col127[11];
                stage2_col127[35] = stage1_col127[11];
                stage2_col127[36] = stage1_col127[11];
                stage2_col127[37] = stage1_col127[11];
                stage2_col127[38] = stage1_col127[11];
                stage2_col127[39] = stage1_col127[11];
                stage2_col127[40] = stage1_col127[11];
                stage2_col127[41] = stage1_col127[11];
                stage2_col127[42] = stage1_col127[11];
                stage2_col127[43] = stage1_col127[11];
                stage2_col127[44] = stage1_col127[11];
                stage2_col127[45] = stage1_col127[11];
                stage2_col127[46] = stage1_col127[11];
                stage2_col127[47] = stage1_col127[11];
                stage2_col127[48] = stage1_col127[11];
                stage2_col127[49] = stage1_col127[11];
            end
        end
    endgenerate

    // Stage 3: Reduction
    fa fa_s2_c4_n0 (
        .a(stage2_col4[0]),
        .b(stage2_col4[1]),
        .c_in(stage2_col4[2]),
        .s(fa_s2_c4_n0_s),
        .c_out(fa_s2_c4_n0_c)
    );

    fa fa_s2_c9_n1 (
        .a(stage2_col9[0]),
        .b(stage2_col9[1]),
        .c_in(stage2_col9[2]),
        .s(fa_s2_c9_n1_s),
        .c_out(fa_s2_c9_n1_c)
    );

    fa fa_s2_c10_n2 (
        .a(stage2_col10[0]),
        .b(stage2_col10[1]),
        .c_in(stage2_col10[2]),
        .s(fa_s2_c10_n2_s),
        .c_out(fa_s2_c10_n2_c)
    );

    fa fa_s2_c11_n3 (
        .a(stage2_col11[0]),
        .b(stage2_col11[1]),
        .c_in(stage2_col11[2]),
        .s(fa_s2_c11_n3_s),
        .c_out(fa_s2_c11_n3_c)
    );

    fa fa_s2_c12_n4 (
        .a(stage2_col12[0]),
        .b(stage2_col12[1]),
        .c_in(stage2_col12[2]),
        .s(fa_s2_c12_n4_s),
        .c_out(fa_s2_c12_n4_c)
    );

    fa fa_s2_c13_n5 (
        .a(stage2_col13[0]),
        .b(stage2_col13[1]),
        .c_in(stage2_col13[2]),
        .s(fa_s2_c13_n5_s),
        .c_out(fa_s2_c13_n5_c)
    );

    fa fa_s2_c14_n6 (
        .a(stage2_col14[0]),
        .b(stage2_col14[1]),
        .c_in(stage2_col14[2]),
        .s(fa_s2_c14_n6_s),
        .c_out(fa_s2_c14_n6_c)
    );

    fa fa_s2_c15_n7 (
        .a(stage2_col15[0]),
        .b(stage2_col15[1]),
        .c_in(stage2_col15[2]),
        .s(fa_s2_c15_n7_s),
        .c_out(fa_s2_c15_n7_c)
    );

    fa fa_s2_c16_n8 (
        .a(stage2_col16[0]),
        .b(stage2_col16[1]),
        .c_in(stage2_col16[2]),
        .s(fa_s2_c16_n8_s),
        .c_out(fa_s2_c16_n8_c)
    );

    fa fa_s2_c17_n9 (
        .a(stage2_col17[0]),
        .b(stage2_col17[1]),
        .c_in(stage2_col17[2]),
        .s(fa_s2_c17_n9_s),
        .c_out(fa_s2_c17_n9_c)
    );

    fa fa_s2_c18_n10 (
        .a(stage2_col18[0]),
        .b(stage2_col18[1]),
        .c_in(stage2_col18[2]),
        .s(fa_s2_c18_n10_s),
        .c_out(fa_s2_c18_n10_c)
    );

    fa fa_s2_c18_n11 (
        .a(stage2_col18[3]),
        .b(stage2_col18[4]),
        .c_in(stage2_col18[5]),
        .s(fa_s2_c18_n11_s),
        .c_out(fa_s2_c18_n11_c)
    );

    fa fa_s2_c19_n12 (
        .a(stage2_col19[0]),
        .b(stage2_col19[1]),
        .c_in(stage2_col19[2]),
        .s(fa_s2_c19_n12_s),
        .c_out(fa_s2_c19_n12_c)
    );

    fa fa_s2_c20_n13 (
        .a(stage2_col20[0]),
        .b(stage2_col20[1]),
        .c_in(stage2_col20[2]),
        .s(fa_s2_c20_n13_s),
        .c_out(fa_s2_c20_n13_c)
    );

    fa fa_s2_c21_n14 (
        .a(stage2_col21[0]),
        .b(stage2_col21[1]),
        .c_in(stage2_col21[2]),
        .s(fa_s2_c21_n14_s),
        .c_out(fa_s2_c21_n14_c)
    );

    fa fa_s2_c22_n15 (
        .a(stage2_col22[0]),
        .b(stage2_col22[1]),
        .c_in(stage2_col22[2]),
        .s(fa_s2_c22_n15_s),
        .c_out(fa_s2_c22_n15_c)
    );

    fa fa_s2_c22_n16 (
        .a(stage2_col22[3]),
        .b(stage2_col22[4]),
        .c_in(stage2_col22[5]),
        .s(fa_s2_c22_n16_s),
        .c_out(fa_s2_c22_n16_c)
    );

    fa fa_s2_c23_n17 (
        .a(stage2_col23[0]),
        .b(stage2_col23[1]),
        .c_in(stage2_col23[2]),
        .s(fa_s2_c23_n17_s),
        .c_out(fa_s2_c23_n17_c)
    );

    fa fa_s2_c23_n18 (
        .a(stage2_col23[3]),
        .b(stage2_col23[4]),
        .c_in(stage2_col23[5]),
        .s(fa_s2_c23_n18_s),
        .c_out(fa_s2_c23_n18_c)
    );

    fa fa_s2_c24_n19 (
        .a(stage2_col24[0]),
        .b(stage2_col24[1]),
        .c_in(stage2_col24[2]),
        .s(fa_s2_c24_n19_s),
        .c_out(fa_s2_c24_n19_c)
    );

    fa fa_s2_c24_n20 (
        .a(stage2_col24[3]),
        .b(stage2_col24[4]),
        .c_in(stage2_col24[5]),
        .s(fa_s2_c24_n20_s),
        .c_out(fa_s2_c24_n20_c)
    );

    fa fa_s2_c25_n21 (
        .a(stage2_col25[0]),
        .b(stage2_col25[1]),
        .c_in(stage2_col25[2]),
        .s(fa_s2_c25_n21_s),
        .c_out(fa_s2_c25_n21_c)
    );

    fa fa_s2_c25_n22 (
        .a(stage2_col25[3]),
        .b(stage2_col25[4]),
        .c_in(stage2_col25[5]),
        .s(fa_s2_c25_n22_s),
        .c_out(fa_s2_c25_n22_c)
    );

    fa fa_s2_c26_n23 (
        .a(stage2_col26[0]),
        .b(stage2_col26[1]),
        .c_in(stage2_col26[2]),
        .s(fa_s2_c26_n23_s),
        .c_out(fa_s2_c26_n23_c)
    );

    fa fa_s2_c26_n24 (
        .a(stage2_col26[3]),
        .b(stage2_col26[4]),
        .c_in(stage2_col26[5]),
        .s(fa_s2_c26_n24_s),
        .c_out(fa_s2_c26_n24_c)
    );

    fa fa_s2_c27_n25 (
        .a(stage2_col27[0]),
        .b(stage2_col27[1]),
        .c_in(stage2_col27[2]),
        .s(fa_s2_c27_n25_s),
        .c_out(fa_s2_c27_n25_c)
    );

    fa fa_s2_c27_n26 (
        .a(stage2_col27[3]),
        .b(stage2_col27[4]),
        .c_in(stage2_col27[5]),
        .s(fa_s2_c27_n26_s),
        .c_out(fa_s2_c27_n26_c)
    );

    fa fa_s2_c28_n27 (
        .a(stage2_col28[0]),
        .b(stage2_col28[1]),
        .c_in(stage2_col28[2]),
        .s(fa_s2_c28_n27_s),
        .c_out(fa_s2_c28_n27_c)
    );

    fa fa_s2_c28_n28 (
        .a(stage2_col28[3]),
        .b(stage2_col28[4]),
        .c_in(stage2_col28[5]),
        .s(fa_s2_c28_n28_s),
        .c_out(fa_s2_c28_n28_c)
    );

    fa fa_s2_c29_n29 (
        .a(stage2_col29[0]),
        .b(stage2_col29[1]),
        .c_in(stage2_col29[2]),
        .s(fa_s2_c29_n29_s),
        .c_out(fa_s2_c29_n29_c)
    );

    fa fa_s2_c29_n30 (
        .a(stage2_col29[3]),
        .b(stage2_col29[4]),
        .c_in(stage2_col29[5]),
        .s(fa_s2_c29_n30_s),
        .c_out(fa_s2_c29_n30_c)
    );

    fa fa_s2_c30_n31 (
        .a(stage2_col30[0]),
        .b(stage2_col30[1]),
        .c_in(stage2_col30[2]),
        .s(fa_s2_c30_n31_s),
        .c_out(fa_s2_c30_n31_c)
    );

    fa fa_s2_c30_n32 (
        .a(stage2_col30[3]),
        .b(stage2_col30[4]),
        .c_in(stage2_col30[5]),
        .s(fa_s2_c30_n32_s),
        .c_out(fa_s2_c30_n32_c)
    );

    fa fa_s2_c31_n33 (
        .a(stage2_col31[0]),
        .b(stage2_col31[1]),
        .c_in(stage2_col31[2]),
        .s(fa_s2_c31_n33_s),
        .c_out(fa_s2_c31_n33_c)
    );

    fa fa_s2_c31_n34 (
        .a(stage2_col31[3]),
        .b(stage2_col31[4]),
        .c_in(stage2_col31[5]),
        .s(fa_s2_c31_n34_s),
        .c_out(fa_s2_c31_n34_c)
    );

    fa fa_s2_c31_n35 (
        .a(stage2_col31[6]),
        .b(stage2_col31[7]),
        .c_in(stage2_col31[8]),
        .s(fa_s2_c31_n35_s),
        .c_out(fa_s2_c31_n35_c)
    );

    fa fa_s2_c32_n36 (
        .a(stage2_col32[0]),
        .b(stage2_col32[1]),
        .c_in(stage2_col32[2]),
        .s(fa_s2_c32_n36_s),
        .c_out(fa_s2_c32_n36_c)
    );

    fa fa_s2_c32_n37 (
        .a(stage2_col32[3]),
        .b(stage2_col32[4]),
        .c_in(stage2_col32[5]),
        .s(fa_s2_c32_n37_s),
        .c_out(fa_s2_c32_n37_c)
    );

    fa fa_s2_c33_n38 (
        .a(stage2_col33[0]),
        .b(stage2_col33[1]),
        .c_in(stage2_col33[2]),
        .s(fa_s2_c33_n38_s),
        .c_out(fa_s2_c33_n38_c)
    );

    fa fa_s2_c33_n39 (
        .a(stage2_col33[3]),
        .b(stage2_col33[4]),
        .c_in(stage2_col33[5]),
        .s(fa_s2_c33_n39_s),
        .c_out(fa_s2_c33_n39_c)
    );

    fa fa_s2_c34_n40 (
        .a(stage2_col34[0]),
        .b(stage2_col34[1]),
        .c_in(stage2_col34[2]),
        .s(fa_s2_c34_n40_s),
        .c_out(fa_s2_c34_n40_c)
    );

    fa fa_s2_c34_n41 (
        .a(stage2_col34[3]),
        .b(stage2_col34[4]),
        .c_in(stage2_col34[5]),
        .s(fa_s2_c34_n41_s),
        .c_out(fa_s2_c34_n41_c)
    );

    fa fa_s2_c35_n42 (
        .a(stage2_col35[0]),
        .b(stage2_col35[1]),
        .c_in(stage2_col35[2]),
        .s(fa_s2_c35_n42_s),
        .c_out(fa_s2_c35_n42_c)
    );

    fa fa_s2_c35_n43 (
        .a(stage2_col35[3]),
        .b(stage2_col35[4]),
        .c_in(stage2_col35[5]),
        .s(fa_s2_c35_n43_s),
        .c_out(fa_s2_c35_n43_c)
    );

    fa fa_s2_c36_n44 (
        .a(stage2_col36[0]),
        .b(stage2_col36[1]),
        .c_in(stage2_col36[2]),
        .s(fa_s2_c36_n44_s),
        .c_out(fa_s2_c36_n44_c)
    );

    fa fa_s2_c36_n45 (
        .a(stage2_col36[3]),
        .b(stage2_col36[4]),
        .c_in(stage2_col36[5]),
        .s(fa_s2_c36_n45_s),
        .c_out(fa_s2_c36_n45_c)
    );

    fa fa_s2_c36_n46 (
        .a(stage2_col36[6]),
        .b(stage2_col36[7]),
        .c_in(stage2_col36[8]),
        .s(fa_s2_c36_n46_s),
        .c_out(fa_s2_c36_n46_c)
    );

    fa fa_s2_c37_n47 (
        .a(stage2_col37[0]),
        .b(stage2_col37[1]),
        .c_in(stage2_col37[2]),
        .s(fa_s2_c37_n47_s),
        .c_out(fa_s2_c37_n47_c)
    );

    fa fa_s2_c37_n48 (
        .a(stage2_col37[3]),
        .b(stage2_col37[4]),
        .c_in(stage2_col37[5]),
        .s(fa_s2_c37_n48_s),
        .c_out(fa_s2_c37_n48_c)
    );

    fa fa_s2_c37_n49 (
        .a(stage2_col37[6]),
        .b(stage2_col37[7]),
        .c_in(stage2_col37[8]),
        .s(fa_s2_c37_n49_s),
        .c_out(fa_s2_c37_n49_c)
    );

    fa fa_s2_c38_n50 (
        .a(stage2_col38[0]),
        .b(stage2_col38[1]),
        .c_in(stage2_col38[2]),
        .s(fa_s2_c38_n50_s),
        .c_out(fa_s2_c38_n50_c)
    );

    fa fa_s2_c38_n51 (
        .a(stage2_col38[3]),
        .b(stage2_col38[4]),
        .c_in(stage2_col38[5]),
        .s(fa_s2_c38_n51_s),
        .c_out(fa_s2_c38_n51_c)
    );

    fa fa_s2_c38_n52 (
        .a(stage2_col38[6]),
        .b(stage2_col38[7]),
        .c_in(stage2_col38[8]),
        .s(fa_s2_c38_n52_s),
        .c_out(fa_s2_c38_n52_c)
    );

    fa fa_s2_c39_n53 (
        .a(stage2_col39[0]),
        .b(stage2_col39[1]),
        .c_in(stage2_col39[2]),
        .s(fa_s2_c39_n53_s),
        .c_out(fa_s2_c39_n53_c)
    );

    fa fa_s2_c39_n54 (
        .a(stage2_col39[3]),
        .b(stage2_col39[4]),
        .c_in(stage2_col39[5]),
        .s(fa_s2_c39_n54_s),
        .c_out(fa_s2_c39_n54_c)
    );

    fa fa_s2_c39_n55 (
        .a(stage2_col39[6]),
        .b(stage2_col39[7]),
        .c_in(stage2_col39[8]),
        .s(fa_s2_c39_n55_s),
        .c_out(fa_s2_c39_n55_c)
    );

    fa fa_s2_c40_n56 (
        .a(stage2_col40[0]),
        .b(stage2_col40[1]),
        .c_in(stage2_col40[2]),
        .s(fa_s2_c40_n56_s),
        .c_out(fa_s2_c40_n56_c)
    );

    fa fa_s2_c40_n57 (
        .a(stage2_col40[3]),
        .b(stage2_col40[4]),
        .c_in(stage2_col40[5]),
        .s(fa_s2_c40_n57_s),
        .c_out(fa_s2_c40_n57_c)
    );

    fa fa_s2_c40_n58 (
        .a(stage2_col40[6]),
        .b(stage2_col40[7]),
        .c_in(stage2_col40[8]),
        .s(fa_s2_c40_n58_s),
        .c_out(fa_s2_c40_n58_c)
    );

    fa fa_s2_c41_n59 (
        .a(stage2_col41[0]),
        .b(stage2_col41[1]),
        .c_in(stage2_col41[2]),
        .s(fa_s2_c41_n59_s),
        .c_out(fa_s2_c41_n59_c)
    );

    fa fa_s2_c41_n60 (
        .a(stage2_col41[3]),
        .b(stage2_col41[4]),
        .c_in(stage2_col41[5]),
        .s(fa_s2_c41_n60_s),
        .c_out(fa_s2_c41_n60_c)
    );

    fa fa_s2_c41_n61 (
        .a(stage2_col41[6]),
        .b(stage2_col41[7]),
        .c_in(stage2_col41[8]),
        .s(fa_s2_c41_n61_s),
        .c_out(fa_s2_c41_n61_c)
    );

    fa fa_s2_c42_n62 (
        .a(stage2_col42[0]),
        .b(stage2_col42[1]),
        .c_in(stage2_col42[2]),
        .s(fa_s2_c42_n62_s),
        .c_out(fa_s2_c42_n62_c)
    );

    fa fa_s2_c42_n63 (
        .a(stage2_col42[3]),
        .b(stage2_col42[4]),
        .c_in(stage2_col42[5]),
        .s(fa_s2_c42_n63_s),
        .c_out(fa_s2_c42_n63_c)
    );

    fa fa_s2_c42_n64 (
        .a(stage2_col42[6]),
        .b(stage2_col42[7]),
        .c_in(stage2_col42[8]),
        .s(fa_s2_c42_n64_s),
        .c_out(fa_s2_c42_n64_c)
    );

    fa fa_s2_c43_n65 (
        .a(stage2_col43[0]),
        .b(stage2_col43[1]),
        .c_in(stage2_col43[2]),
        .s(fa_s2_c43_n65_s),
        .c_out(fa_s2_c43_n65_c)
    );

    fa fa_s2_c43_n66 (
        .a(stage2_col43[3]),
        .b(stage2_col43[4]),
        .c_in(stage2_col43[5]),
        .s(fa_s2_c43_n66_s),
        .c_out(fa_s2_c43_n66_c)
    );

    fa fa_s2_c43_n67 (
        .a(stage2_col43[6]),
        .b(stage2_col43[7]),
        .c_in(stage2_col43[8]),
        .s(fa_s2_c43_n67_s),
        .c_out(fa_s2_c43_n67_c)
    );

    fa fa_s2_c44_n68 (
        .a(stage2_col44[0]),
        .b(stage2_col44[1]),
        .c_in(stage2_col44[2]),
        .s(fa_s2_c44_n68_s),
        .c_out(fa_s2_c44_n68_c)
    );

    fa fa_s2_c44_n69 (
        .a(stage2_col44[3]),
        .b(stage2_col44[4]),
        .c_in(stage2_col44[5]),
        .s(fa_s2_c44_n69_s),
        .c_out(fa_s2_c44_n69_c)
    );

    fa fa_s2_c44_n70 (
        .a(stage2_col44[6]),
        .b(stage2_col44[7]),
        .c_in(stage2_col44[8]),
        .s(fa_s2_c44_n70_s),
        .c_out(fa_s2_c44_n70_c)
    );

    fa fa_s2_c45_n71 (
        .a(stage2_col45[0]),
        .b(stage2_col45[1]),
        .c_in(stage2_col45[2]),
        .s(fa_s2_c45_n71_s),
        .c_out(fa_s2_c45_n71_c)
    );

    fa fa_s2_c45_n72 (
        .a(stage2_col45[3]),
        .b(stage2_col45[4]),
        .c_in(stage2_col45[5]),
        .s(fa_s2_c45_n72_s),
        .c_out(fa_s2_c45_n72_c)
    );

    fa fa_s2_c45_n73 (
        .a(stage2_col45[6]),
        .b(stage2_col45[7]),
        .c_in(stage2_col45[8]),
        .s(fa_s2_c45_n73_s),
        .c_out(fa_s2_c45_n73_c)
    );

    fa fa_s2_c45_n74 (
        .a(stage2_col45[9]),
        .b(stage2_col45[10]),
        .c_in(stage2_col45[11]),
        .s(fa_s2_c45_n74_s),
        .c_out(fa_s2_c45_n74_c)
    );

    fa fa_s2_c46_n75 (
        .a(stage2_col46[0]),
        .b(stage2_col46[1]),
        .c_in(stage2_col46[2]),
        .s(fa_s2_c46_n75_s),
        .c_out(fa_s2_c46_n75_c)
    );

    fa fa_s2_c46_n76 (
        .a(stage2_col46[3]),
        .b(stage2_col46[4]),
        .c_in(stage2_col46[5]),
        .s(fa_s2_c46_n76_s),
        .c_out(fa_s2_c46_n76_c)
    );

    fa fa_s2_c46_n77 (
        .a(stage2_col46[6]),
        .b(stage2_col46[7]),
        .c_in(stage2_col46[8]),
        .s(fa_s2_c46_n77_s),
        .c_out(fa_s2_c46_n77_c)
    );

    fa fa_s2_c47_n78 (
        .a(stage2_col47[0]),
        .b(stage2_col47[1]),
        .c_in(stage2_col47[2]),
        .s(fa_s2_c47_n78_s),
        .c_out(fa_s2_c47_n78_c)
    );

    fa fa_s2_c47_n79 (
        .a(stage2_col47[3]),
        .b(stage2_col47[4]),
        .c_in(stage2_col47[5]),
        .s(fa_s2_c47_n79_s),
        .c_out(fa_s2_c47_n79_c)
    );

    fa fa_s2_c47_n80 (
        .a(stage2_col47[6]),
        .b(stage2_col47[7]),
        .c_in(stage2_col47[8]),
        .s(fa_s2_c47_n80_s),
        .c_out(fa_s2_c47_n80_c)
    );

    fa fa_s2_c48_n81 (
        .a(stage2_col48[0]),
        .b(stage2_col48[1]),
        .c_in(stage2_col48[2]),
        .s(fa_s2_c48_n81_s),
        .c_out(fa_s2_c48_n81_c)
    );

    fa fa_s2_c48_n82 (
        .a(stage2_col48[3]),
        .b(stage2_col48[4]),
        .c_in(stage2_col48[5]),
        .s(fa_s2_c48_n82_s),
        .c_out(fa_s2_c48_n82_c)
    );

    fa fa_s2_c48_n83 (
        .a(stage2_col48[6]),
        .b(stage2_col48[7]),
        .c_in(stage2_col48[8]),
        .s(fa_s2_c48_n83_s),
        .c_out(fa_s2_c48_n83_c)
    );

    fa fa_s2_c49_n84 (
        .a(stage2_col49[0]),
        .b(stage2_col49[1]),
        .c_in(stage2_col49[2]),
        .s(fa_s2_c49_n84_s),
        .c_out(fa_s2_c49_n84_c)
    );

    fa fa_s2_c49_n85 (
        .a(stage2_col49[3]),
        .b(stage2_col49[4]),
        .c_in(stage2_col49[5]),
        .s(fa_s2_c49_n85_s),
        .c_out(fa_s2_c49_n85_c)
    );

    fa fa_s2_c49_n86 (
        .a(stage2_col49[6]),
        .b(stage2_col49[7]),
        .c_in(stage2_col49[8]),
        .s(fa_s2_c49_n86_s),
        .c_out(fa_s2_c49_n86_c)
    );

    fa fa_s2_c49_n87 (
        .a(stage2_col49[9]),
        .b(stage2_col49[10]),
        .c_in(stage2_col49[11]),
        .s(fa_s2_c49_n87_s),
        .c_out(fa_s2_c49_n87_c)
    );

    fa fa_s2_c50_n88 (
        .a(stage2_col50[0]),
        .b(stage2_col50[1]),
        .c_in(stage2_col50[2]),
        .s(fa_s2_c50_n88_s),
        .c_out(fa_s2_c50_n88_c)
    );

    fa fa_s2_c50_n89 (
        .a(stage2_col50[3]),
        .b(stage2_col50[4]),
        .c_in(stage2_col50[5]),
        .s(fa_s2_c50_n89_s),
        .c_out(fa_s2_c50_n89_c)
    );

    fa fa_s2_c50_n90 (
        .a(stage2_col50[6]),
        .b(stage2_col50[7]),
        .c_in(stage2_col50[8]),
        .s(fa_s2_c50_n90_s),
        .c_out(fa_s2_c50_n90_c)
    );

    fa fa_s2_c50_n91 (
        .a(stage2_col50[9]),
        .b(stage2_col50[10]),
        .c_in(stage2_col50[11]),
        .s(fa_s2_c50_n91_s),
        .c_out(fa_s2_c50_n91_c)
    );

    fa fa_s2_c51_n92 (
        .a(stage2_col51[0]),
        .b(stage2_col51[1]),
        .c_in(stage2_col51[2]),
        .s(fa_s2_c51_n92_s),
        .c_out(fa_s2_c51_n92_c)
    );

    fa fa_s2_c51_n93 (
        .a(stage2_col51[3]),
        .b(stage2_col51[4]),
        .c_in(stage2_col51[5]),
        .s(fa_s2_c51_n93_s),
        .c_out(fa_s2_c51_n93_c)
    );

    fa fa_s2_c51_n94 (
        .a(stage2_col51[6]),
        .b(stage2_col51[7]),
        .c_in(stage2_col51[8]),
        .s(fa_s2_c51_n94_s),
        .c_out(fa_s2_c51_n94_c)
    );

    fa fa_s2_c51_n95 (
        .a(stage2_col51[9]),
        .b(stage2_col51[10]),
        .c_in(stage2_col51[11]),
        .s(fa_s2_c51_n95_s),
        .c_out(fa_s2_c51_n95_c)
    );

    fa fa_s2_c52_n96 (
        .a(stage2_col52[0]),
        .b(stage2_col52[1]),
        .c_in(stage2_col52[2]),
        .s(fa_s2_c52_n96_s),
        .c_out(fa_s2_c52_n96_c)
    );

    fa fa_s2_c52_n97 (
        .a(stage2_col52[3]),
        .b(stage2_col52[4]),
        .c_in(stage2_col52[5]),
        .s(fa_s2_c52_n97_s),
        .c_out(fa_s2_c52_n97_c)
    );

    fa fa_s2_c52_n98 (
        .a(stage2_col52[6]),
        .b(stage2_col52[7]),
        .c_in(stage2_col52[8]),
        .s(fa_s2_c52_n98_s),
        .c_out(fa_s2_c52_n98_c)
    );

    fa fa_s2_c52_n99 (
        .a(stage2_col52[9]),
        .b(stage2_col52[10]),
        .c_in(stage2_col52[11]),
        .s(fa_s2_c52_n99_s),
        .c_out(fa_s2_c52_n99_c)
    );

    fa fa_s2_c53_n100 (
        .a(stage2_col53[0]),
        .b(stage2_col53[1]),
        .c_in(stage2_col53[2]),
        .s(fa_s2_c53_n100_s),
        .c_out(fa_s2_c53_n100_c)
    );

    fa fa_s2_c53_n101 (
        .a(stage2_col53[3]),
        .b(stage2_col53[4]),
        .c_in(stage2_col53[5]),
        .s(fa_s2_c53_n101_s),
        .c_out(fa_s2_c53_n101_c)
    );

    fa fa_s2_c53_n102 (
        .a(stage2_col53[6]),
        .b(stage2_col53[7]),
        .c_in(stage2_col53[8]),
        .s(fa_s2_c53_n102_s),
        .c_out(fa_s2_c53_n102_c)
    );

    fa fa_s2_c53_n103 (
        .a(stage2_col53[9]),
        .b(stage2_col53[10]),
        .c_in(stage2_col53[11]),
        .s(fa_s2_c53_n103_s),
        .c_out(fa_s2_c53_n103_c)
    );

    fa fa_s2_c54_n104 (
        .a(stage2_col54[0]),
        .b(stage2_col54[1]),
        .c_in(stage2_col54[2]),
        .s(fa_s2_c54_n104_s),
        .c_out(fa_s2_c54_n104_c)
    );

    fa fa_s2_c54_n105 (
        .a(stage2_col54[3]),
        .b(stage2_col54[4]),
        .c_in(stage2_col54[5]),
        .s(fa_s2_c54_n105_s),
        .c_out(fa_s2_c54_n105_c)
    );

    fa fa_s2_c54_n106 (
        .a(stage2_col54[6]),
        .b(stage2_col54[7]),
        .c_in(stage2_col54[8]),
        .s(fa_s2_c54_n106_s),
        .c_out(fa_s2_c54_n106_c)
    );

    fa fa_s2_c54_n107 (
        .a(stage2_col54[9]),
        .b(stage2_col54[10]),
        .c_in(stage2_col54[11]),
        .s(fa_s2_c54_n107_s),
        .c_out(fa_s2_c54_n107_c)
    );

    fa fa_s2_c55_n108 (
        .a(stage2_col55[0]),
        .b(stage2_col55[1]),
        .c_in(stage2_col55[2]),
        .s(fa_s2_c55_n108_s),
        .c_out(fa_s2_c55_n108_c)
    );

    fa fa_s2_c55_n109 (
        .a(stage2_col55[3]),
        .b(stage2_col55[4]),
        .c_in(stage2_col55[5]),
        .s(fa_s2_c55_n109_s),
        .c_out(fa_s2_c55_n109_c)
    );

    fa fa_s2_c55_n110 (
        .a(stage2_col55[6]),
        .b(stage2_col55[7]),
        .c_in(stage2_col55[8]),
        .s(fa_s2_c55_n110_s),
        .c_out(fa_s2_c55_n110_c)
    );

    fa fa_s2_c55_n111 (
        .a(stage2_col55[9]),
        .b(stage2_col55[10]),
        .c_in(stage2_col55[11]),
        .s(fa_s2_c55_n111_s),
        .c_out(fa_s2_c55_n111_c)
    );

    fa fa_s2_c56_n112 (
        .a(stage2_col56[0]),
        .b(stage2_col56[1]),
        .c_in(stage2_col56[2]),
        .s(fa_s2_c56_n112_s),
        .c_out(fa_s2_c56_n112_c)
    );

    fa fa_s2_c56_n113 (
        .a(stage2_col56[3]),
        .b(stage2_col56[4]),
        .c_in(stage2_col56[5]),
        .s(fa_s2_c56_n113_s),
        .c_out(fa_s2_c56_n113_c)
    );

    fa fa_s2_c56_n114 (
        .a(stage2_col56[6]),
        .b(stage2_col56[7]),
        .c_in(stage2_col56[8]),
        .s(fa_s2_c56_n114_s),
        .c_out(fa_s2_c56_n114_c)
    );

    fa fa_s2_c56_n115 (
        .a(stage2_col56[9]),
        .b(stage2_col56[10]),
        .c_in(stage2_col56[11]),
        .s(fa_s2_c56_n115_s),
        .c_out(fa_s2_c56_n115_c)
    );

    fa fa_s2_c57_n116 (
        .a(stage2_col57[0]),
        .b(stage2_col57[1]),
        .c_in(stage2_col57[2]),
        .s(fa_s2_c57_n116_s),
        .c_out(fa_s2_c57_n116_c)
    );

    fa fa_s2_c57_n117 (
        .a(stage2_col57[3]),
        .b(stage2_col57[4]),
        .c_in(stage2_col57[5]),
        .s(fa_s2_c57_n117_s),
        .c_out(fa_s2_c57_n117_c)
    );

    fa fa_s2_c57_n118 (
        .a(stage2_col57[6]),
        .b(stage2_col57[7]),
        .c_in(stage2_col57[8]),
        .s(fa_s2_c57_n118_s),
        .c_out(fa_s2_c57_n118_c)
    );

    fa fa_s2_c57_n119 (
        .a(stage2_col57[9]),
        .b(stage2_col57[10]),
        .c_in(stage2_col57[11]),
        .s(fa_s2_c57_n119_s),
        .c_out(fa_s2_c57_n119_c)
    );

    fa fa_s2_c58_n120 (
        .a(stage2_col58[0]),
        .b(stage2_col58[1]),
        .c_in(stage2_col58[2]),
        .s(fa_s2_c58_n120_s),
        .c_out(fa_s2_c58_n120_c)
    );

    fa fa_s2_c58_n121 (
        .a(stage2_col58[3]),
        .b(stage2_col58[4]),
        .c_in(stage2_col58[5]),
        .s(fa_s2_c58_n121_s),
        .c_out(fa_s2_c58_n121_c)
    );

    fa fa_s2_c58_n122 (
        .a(stage2_col58[6]),
        .b(stage2_col58[7]),
        .c_in(stage2_col58[8]),
        .s(fa_s2_c58_n122_s),
        .c_out(fa_s2_c58_n122_c)
    );

    fa fa_s2_c58_n123 (
        .a(stage2_col58[9]),
        .b(stage2_col58[10]),
        .c_in(stage2_col58[11]),
        .s(fa_s2_c58_n123_s),
        .c_out(fa_s2_c58_n123_c)
    );

    fa fa_s2_c58_n124 (
        .a(stage2_col58[12]),
        .b(stage2_col58[13]),
        .c_in(stage2_col58[14]),
        .s(fa_s2_c58_n124_s),
        .c_out(fa_s2_c58_n124_c)
    );

    fa fa_s2_c59_n125 (
        .a(stage2_col59[0]),
        .b(stage2_col59[1]),
        .c_in(stage2_col59[2]),
        .s(fa_s2_c59_n125_s),
        .c_out(fa_s2_c59_n125_c)
    );

    fa fa_s2_c59_n126 (
        .a(stage2_col59[3]),
        .b(stage2_col59[4]),
        .c_in(stage2_col59[5]),
        .s(fa_s2_c59_n126_s),
        .c_out(fa_s2_c59_n126_c)
    );

    fa fa_s2_c59_n127 (
        .a(stage2_col59[6]),
        .b(stage2_col59[7]),
        .c_in(stage2_col59[8]),
        .s(fa_s2_c59_n127_s),
        .c_out(fa_s2_c59_n127_c)
    );

    fa fa_s2_c59_n128 (
        .a(stage2_col59[9]),
        .b(stage2_col59[10]),
        .c_in(stage2_col59[11]),
        .s(fa_s2_c59_n128_s),
        .c_out(fa_s2_c59_n128_c)
    );

    fa fa_s2_c60_n129 (
        .a(stage2_col60[0]),
        .b(stage2_col60[1]),
        .c_in(stage2_col60[2]),
        .s(fa_s2_c60_n129_s),
        .c_out(fa_s2_c60_n129_c)
    );

    fa fa_s2_c60_n130 (
        .a(stage2_col60[3]),
        .b(stage2_col60[4]),
        .c_in(stage2_col60[5]),
        .s(fa_s2_c60_n130_s),
        .c_out(fa_s2_c60_n130_c)
    );

    fa fa_s2_c60_n131 (
        .a(stage2_col60[6]),
        .b(stage2_col60[7]),
        .c_in(stage2_col60[8]),
        .s(fa_s2_c60_n131_s),
        .c_out(fa_s2_c60_n131_c)
    );

    fa fa_s2_c60_n132 (
        .a(stage2_col60[9]),
        .b(stage2_col60[10]),
        .c_in(stage2_col60[11]),
        .s(fa_s2_c60_n132_s),
        .c_out(fa_s2_c60_n132_c)
    );

    fa fa_s2_c61_n133 (
        .a(stage2_col61[0]),
        .b(stage2_col61[1]),
        .c_in(stage2_col61[2]),
        .s(fa_s2_c61_n133_s),
        .c_out(fa_s2_c61_n133_c)
    );

    fa fa_s2_c61_n134 (
        .a(stage2_col61[3]),
        .b(stage2_col61[4]),
        .c_in(stage2_col61[5]),
        .s(fa_s2_c61_n134_s),
        .c_out(fa_s2_c61_n134_c)
    );

    fa fa_s2_c61_n135 (
        .a(stage2_col61[6]),
        .b(stage2_col61[7]),
        .c_in(stage2_col61[8]),
        .s(fa_s2_c61_n135_s),
        .c_out(fa_s2_c61_n135_c)
    );

    fa fa_s2_c61_n136 (
        .a(stage2_col61[9]),
        .b(stage2_col61[10]),
        .c_in(stage2_col61[11]),
        .s(fa_s2_c61_n136_s),
        .c_out(fa_s2_c61_n136_c)
    );

    fa fa_s2_c62_n137 (
        .a(stage2_col62[0]),
        .b(stage2_col62[1]),
        .c_in(stage2_col62[2]),
        .s(fa_s2_c62_n137_s),
        .c_out(fa_s2_c62_n137_c)
    );

    fa fa_s2_c62_n138 (
        .a(stage2_col62[3]),
        .b(stage2_col62[4]),
        .c_in(stage2_col62[5]),
        .s(fa_s2_c62_n138_s),
        .c_out(fa_s2_c62_n138_c)
    );

    fa fa_s2_c62_n139 (
        .a(stage2_col62[6]),
        .b(stage2_col62[7]),
        .c_in(stage2_col62[8]),
        .s(fa_s2_c62_n139_s),
        .c_out(fa_s2_c62_n139_c)
    );

    fa fa_s2_c62_n140 (
        .a(stage2_col62[9]),
        .b(stage2_col62[10]),
        .c_in(stage2_col62[11]),
        .s(fa_s2_c62_n140_s),
        .c_out(fa_s2_c62_n140_c)
    );

    fa fa_s2_c63_n141 (
        .a(stage2_col63[0]),
        .b(stage2_col63[1]),
        .c_in(stage2_col63[2]),
        .s(fa_s2_c63_n141_s),
        .c_out(fa_s2_c63_n141_c)
    );

    fa fa_s2_c63_n142 (
        .a(stage2_col63[3]),
        .b(stage2_col63[4]),
        .c_in(stage2_col63[5]),
        .s(fa_s2_c63_n142_s),
        .c_out(fa_s2_c63_n142_c)
    );

    fa fa_s2_c63_n143 (
        .a(stage2_col63[6]),
        .b(stage2_col63[7]),
        .c_in(stage2_col63[8]),
        .s(fa_s2_c63_n143_s),
        .c_out(fa_s2_c63_n143_c)
    );

    fa fa_s2_c63_n144 (
        .a(stage2_col63[9]),
        .b(stage2_col63[10]),
        .c_in(stage2_col63[11]),
        .s(fa_s2_c63_n144_s),
        .c_out(fa_s2_c63_n144_c)
    );

    fa fa_s2_c63_n145 (
        .a(stage2_col63[12]),
        .b(stage2_col63[13]),
        .c_in(stage2_col63[14]),
        .s(fa_s2_c63_n145_s),
        .c_out(fa_s2_c63_n145_c)
    );

    fa fa_s2_c64_n146 (
        .a(stage2_col64[0]),
        .b(stage2_col64[1]),
        .c_in(stage2_col64[2]),
        .s(fa_s2_c64_n146_s),
        .c_out(fa_s2_c64_n146_c)
    );

    fa fa_s2_c64_n147 (
        .a(stage2_col64[3]),
        .b(stage2_col64[4]),
        .c_in(stage2_col64[5]),
        .s(fa_s2_c64_n147_s),
        .c_out(fa_s2_c64_n147_c)
    );

    fa fa_s2_c64_n148 (
        .a(stage2_col64[6]),
        .b(stage2_col64[7]),
        .c_in(stage2_col64[8]),
        .s(fa_s2_c64_n148_s),
        .c_out(fa_s2_c64_n148_c)
    );

    fa fa_s2_c64_n149 (
        .a(stage2_col64[9]),
        .b(stage2_col64[10]),
        .c_in(stage2_col64[11]),
        .s(fa_s2_c64_n149_s),
        .c_out(fa_s2_c64_n149_c)
    );

    fa fa_s2_c65_n150 (
        .a(stage2_col65[0]),
        .b(stage2_col65[1]),
        .c_in(stage2_col65[2]),
        .s(fa_s2_c65_n150_s),
        .c_out(fa_s2_c65_n150_c)
    );

    fa fa_s2_c65_n151 (
        .a(stage2_col65[3]),
        .b(stage2_col65[4]),
        .c_in(stage2_col65[5]),
        .s(fa_s2_c65_n151_s),
        .c_out(fa_s2_c65_n151_c)
    );

    fa fa_s2_c65_n152 (
        .a(stage2_col65[6]),
        .b(stage2_col65[7]),
        .c_in(stage2_col65[8]),
        .s(fa_s2_c65_n152_s),
        .c_out(fa_s2_c65_n152_c)
    );

    fa fa_s2_c65_n153 (
        .a(stage2_col65[9]),
        .b(stage2_col65[10]),
        .c_in(stage2_col65[11]),
        .s(fa_s2_c65_n153_s),
        .c_out(fa_s2_c65_n153_c)
    );

    fa fa_s2_c65_n154 (
        .a(stage2_col65[12]),
        .b(stage2_col65[13]),
        .c_in(stage2_col65[14]),
        .s(fa_s2_c65_n154_s),
        .c_out(fa_s2_c65_n154_c)
    );

    fa fa_s2_c66_n155 (
        .a(stage2_col66[0]),
        .b(stage2_col66[1]),
        .c_in(stage2_col66[2]),
        .s(fa_s2_c66_n155_s),
        .c_out(fa_s2_c66_n155_c)
    );

    fa fa_s2_c66_n156 (
        .a(stage2_col66[3]),
        .b(stage2_col66[4]),
        .c_in(stage2_col66[5]),
        .s(fa_s2_c66_n156_s),
        .c_out(fa_s2_c66_n156_c)
    );

    fa fa_s2_c66_n157 (
        .a(stage2_col66[6]),
        .b(stage2_col66[7]),
        .c_in(stage2_col66[8]),
        .s(fa_s2_c66_n157_s),
        .c_out(fa_s2_c66_n157_c)
    );

    fa fa_s2_c66_n158 (
        .a(stage2_col66[9]),
        .b(stage2_col66[10]),
        .c_in(stage2_col66[11]),
        .s(fa_s2_c66_n158_s),
        .c_out(fa_s2_c66_n158_c)
    );

    fa fa_s2_c67_n159 (
        .a(stage2_col67[0]),
        .b(stage2_col67[1]),
        .c_in(stage2_col67[2]),
        .s(fa_s2_c67_n159_s),
        .c_out(fa_s2_c67_n159_c)
    );

    fa fa_s2_c67_n160 (
        .a(stage2_col67[3]),
        .b(stage2_col67[4]),
        .c_in(stage2_col67[5]),
        .s(fa_s2_c67_n160_s),
        .c_out(fa_s2_c67_n160_c)
    );

    fa fa_s2_c67_n161 (
        .a(stage2_col67[6]),
        .b(stage2_col67[7]),
        .c_in(stage2_col67[8]),
        .s(fa_s2_c67_n161_s),
        .c_out(fa_s2_c67_n161_c)
    );

    fa fa_s2_c67_n162 (
        .a(stage2_col67[9]),
        .b(stage2_col67[10]),
        .c_in(stage2_col67[11]),
        .s(fa_s2_c67_n162_s),
        .c_out(fa_s2_c67_n162_c)
    );

    fa fa_s2_c67_n163 (
        .a(stage2_col67[12]),
        .b(stage2_col67[13]),
        .c_in(stage2_col67[14]),
        .s(fa_s2_c67_n163_s),
        .c_out(fa_s2_c67_n163_c)
    );

    fa fa_s2_c68_n164 (
        .a(stage2_col68[0]),
        .b(stage2_col68[1]),
        .c_in(stage2_col68[2]),
        .s(fa_s2_c68_n164_s),
        .c_out(fa_s2_c68_n164_c)
    );

    fa fa_s2_c68_n165 (
        .a(stage2_col68[3]),
        .b(stage2_col68[4]),
        .c_in(stage2_col68[5]),
        .s(fa_s2_c68_n165_s),
        .c_out(fa_s2_c68_n165_c)
    );

    fa fa_s2_c68_n166 (
        .a(stage2_col68[6]),
        .b(stage2_col68[7]),
        .c_in(stage2_col68[8]),
        .s(fa_s2_c68_n166_s),
        .c_out(fa_s2_c68_n166_c)
    );

    fa fa_s2_c68_n167 (
        .a(stage2_col68[9]),
        .b(stage2_col68[10]),
        .c_in(stage2_col68[11]),
        .s(fa_s2_c68_n167_s),
        .c_out(fa_s2_c68_n167_c)
    );

    fa fa_s2_c69_n168 (
        .a(stage2_col69[0]),
        .b(stage2_col69[1]),
        .c_in(stage2_col69[2]),
        .s(fa_s2_c69_n168_s),
        .c_out(fa_s2_c69_n168_c)
    );

    fa fa_s2_c69_n169 (
        .a(stage2_col69[3]),
        .b(stage2_col69[4]),
        .c_in(stage2_col69[5]),
        .s(fa_s2_c69_n169_s),
        .c_out(fa_s2_c69_n169_c)
    );

    fa fa_s2_c69_n170 (
        .a(stage2_col69[6]),
        .b(stage2_col69[7]),
        .c_in(stage2_col69[8]),
        .s(fa_s2_c69_n170_s),
        .c_out(fa_s2_c69_n170_c)
    );

    fa fa_s2_c69_n171 (
        .a(stage2_col69[9]),
        .b(stage2_col69[10]),
        .c_in(stage2_col69[11]),
        .s(fa_s2_c69_n171_s),
        .c_out(fa_s2_c69_n171_c)
    );

    fa fa_s2_c69_n172 (
        .a(stage2_col69[12]),
        .b(stage2_col69[13]),
        .c_in(stage2_col69[14]),
        .s(fa_s2_c69_n172_s),
        .c_out(fa_s2_c69_n172_c)
    );

    fa fa_s2_c70_n173 (
        .a(stage2_col70[0]),
        .b(stage2_col70[1]),
        .c_in(stage2_col70[2]),
        .s(fa_s2_c70_n173_s),
        .c_out(fa_s2_c70_n173_c)
    );

    fa fa_s2_c70_n174 (
        .a(stage2_col70[3]),
        .b(stage2_col70[4]),
        .c_in(stage2_col70[5]),
        .s(fa_s2_c70_n174_s),
        .c_out(fa_s2_c70_n174_c)
    );

    fa fa_s2_c70_n175 (
        .a(stage2_col70[6]),
        .b(stage2_col70[7]),
        .c_in(stage2_col70[8]),
        .s(fa_s2_c70_n175_s),
        .c_out(fa_s2_c70_n175_c)
    );

    fa fa_s2_c70_n176 (
        .a(stage2_col70[9]),
        .b(stage2_col70[10]),
        .c_in(stage2_col70[11]),
        .s(fa_s2_c70_n176_s),
        .c_out(fa_s2_c70_n176_c)
    );

    fa fa_s2_c71_n177 (
        .a(stage2_col71[0]),
        .b(stage2_col71[1]),
        .c_in(stage2_col71[2]),
        .s(fa_s2_c71_n177_s),
        .c_out(fa_s2_c71_n177_c)
    );

    fa fa_s2_c71_n178 (
        .a(stage2_col71[3]),
        .b(stage2_col71[4]),
        .c_in(stage2_col71[5]),
        .s(fa_s2_c71_n178_s),
        .c_out(fa_s2_c71_n178_c)
    );

    fa fa_s2_c71_n179 (
        .a(stage2_col71[6]),
        .b(stage2_col71[7]),
        .c_in(stage2_col71[8]),
        .s(fa_s2_c71_n179_s),
        .c_out(fa_s2_c71_n179_c)
    );

    fa fa_s2_c71_n180 (
        .a(stage2_col71[9]),
        .b(stage2_col71[10]),
        .c_in(stage2_col71[11]),
        .s(fa_s2_c71_n180_s),
        .c_out(fa_s2_c71_n180_c)
    );

    fa fa_s2_c71_n181 (
        .a(stage2_col71[12]),
        .b(stage2_col71[13]),
        .c_in(stage2_col71[14]),
        .s(fa_s2_c71_n181_s),
        .c_out(fa_s2_c71_n181_c)
    );

    fa fa_s2_c72_n182 (
        .a(stage2_col72[0]),
        .b(stage2_col72[1]),
        .c_in(stage2_col72[2]),
        .s(fa_s2_c72_n182_s),
        .c_out(fa_s2_c72_n182_c)
    );

    fa fa_s2_c72_n183 (
        .a(stage2_col72[3]),
        .b(stage2_col72[4]),
        .c_in(stage2_col72[5]),
        .s(fa_s2_c72_n183_s),
        .c_out(fa_s2_c72_n183_c)
    );

    fa fa_s2_c72_n184 (
        .a(stage2_col72[6]),
        .b(stage2_col72[7]),
        .c_in(stage2_col72[8]),
        .s(fa_s2_c72_n184_s),
        .c_out(fa_s2_c72_n184_c)
    );

    fa fa_s2_c72_n185 (
        .a(stage2_col72[9]),
        .b(stage2_col72[10]),
        .c_in(stage2_col72[11]),
        .s(fa_s2_c72_n185_s),
        .c_out(fa_s2_c72_n185_c)
    );

    fa fa_s2_c73_n186 (
        .a(stage2_col73[0]),
        .b(stage2_col73[1]),
        .c_in(stage2_col73[2]),
        .s(fa_s2_c73_n186_s),
        .c_out(fa_s2_c73_n186_c)
    );

    fa fa_s2_c73_n187 (
        .a(stage2_col73[3]),
        .b(stage2_col73[4]),
        .c_in(stage2_col73[5]),
        .s(fa_s2_c73_n187_s),
        .c_out(fa_s2_c73_n187_c)
    );

    fa fa_s2_c73_n188 (
        .a(stage2_col73[6]),
        .b(stage2_col73[7]),
        .c_in(stage2_col73[8]),
        .s(fa_s2_c73_n188_s),
        .c_out(fa_s2_c73_n188_c)
    );

    fa fa_s2_c73_n189 (
        .a(stage2_col73[9]),
        .b(stage2_col73[10]),
        .c_in(stage2_col73[11]),
        .s(fa_s2_c73_n189_s),
        .c_out(fa_s2_c73_n189_c)
    );

    fa fa_s2_c73_n190 (
        .a(stage2_col73[12]),
        .b(stage2_col73[13]),
        .c_in(stage2_col73[14]),
        .s(fa_s2_c73_n190_s),
        .c_out(fa_s2_c73_n190_c)
    );

    fa fa_s2_c74_n191 (
        .a(stage2_col74[0]),
        .b(stage2_col74[1]),
        .c_in(stage2_col74[2]),
        .s(fa_s2_c74_n191_s),
        .c_out(fa_s2_c74_n191_c)
    );

    fa fa_s2_c74_n192 (
        .a(stage2_col74[3]),
        .b(stage2_col74[4]),
        .c_in(stage2_col74[5]),
        .s(fa_s2_c74_n192_s),
        .c_out(fa_s2_c74_n192_c)
    );

    fa fa_s2_c74_n193 (
        .a(stage2_col74[6]),
        .b(stage2_col74[7]),
        .c_in(stage2_col74[8]),
        .s(fa_s2_c74_n193_s),
        .c_out(fa_s2_c74_n193_c)
    );

    fa fa_s2_c74_n194 (
        .a(stage2_col74[9]),
        .b(stage2_col74[10]),
        .c_in(stage2_col74[11]),
        .s(fa_s2_c74_n194_s),
        .c_out(fa_s2_c74_n194_c)
    );

    fa fa_s2_c75_n195 (
        .a(stage2_col75[0]),
        .b(stage2_col75[1]),
        .c_in(stage2_col75[2]),
        .s(fa_s2_c75_n195_s),
        .c_out(fa_s2_c75_n195_c)
    );

    fa fa_s2_c75_n196 (
        .a(stage2_col75[3]),
        .b(stage2_col75[4]),
        .c_in(stage2_col75[5]),
        .s(fa_s2_c75_n196_s),
        .c_out(fa_s2_c75_n196_c)
    );

    fa fa_s2_c75_n197 (
        .a(stage2_col75[6]),
        .b(stage2_col75[7]),
        .c_in(stage2_col75[8]),
        .s(fa_s2_c75_n197_s),
        .c_out(fa_s2_c75_n197_c)
    );

    fa fa_s2_c75_n198 (
        .a(stage2_col75[9]),
        .b(stage2_col75[10]),
        .c_in(stage2_col75[11]),
        .s(fa_s2_c75_n198_s),
        .c_out(fa_s2_c75_n198_c)
    );

    fa fa_s2_c75_n199 (
        .a(stage2_col75[12]),
        .b(stage2_col75[13]),
        .c_in(stage2_col75[14]),
        .s(fa_s2_c75_n199_s),
        .c_out(fa_s2_c75_n199_c)
    );

    fa fa_s2_c76_n200 (
        .a(stage2_col76[0]),
        .b(stage2_col76[1]),
        .c_in(stage2_col76[2]),
        .s(fa_s2_c76_n200_s),
        .c_out(fa_s2_c76_n200_c)
    );

    fa fa_s2_c76_n201 (
        .a(stage2_col76[3]),
        .b(stage2_col76[4]),
        .c_in(stage2_col76[5]),
        .s(fa_s2_c76_n201_s),
        .c_out(fa_s2_c76_n201_c)
    );

    fa fa_s2_c76_n202 (
        .a(stage2_col76[6]),
        .b(stage2_col76[7]),
        .c_in(stage2_col76[8]),
        .s(fa_s2_c76_n202_s),
        .c_out(fa_s2_c76_n202_c)
    );

    fa fa_s2_c76_n203 (
        .a(stage2_col76[9]),
        .b(stage2_col76[10]),
        .c_in(stage2_col76[11]),
        .s(fa_s2_c76_n203_s),
        .c_out(fa_s2_c76_n203_c)
    );

    fa fa_s2_c77_n204 (
        .a(stage2_col77[0]),
        .b(stage2_col77[1]),
        .c_in(stage2_col77[2]),
        .s(fa_s2_c77_n204_s),
        .c_out(fa_s2_c77_n204_c)
    );

    fa fa_s2_c77_n205 (
        .a(stage2_col77[3]),
        .b(stage2_col77[4]),
        .c_in(stage2_col77[5]),
        .s(fa_s2_c77_n205_s),
        .c_out(fa_s2_c77_n205_c)
    );

    fa fa_s2_c77_n206 (
        .a(stage2_col77[6]),
        .b(stage2_col77[7]),
        .c_in(stage2_col77[8]),
        .s(fa_s2_c77_n206_s),
        .c_out(fa_s2_c77_n206_c)
    );

    fa fa_s2_c77_n207 (
        .a(stage2_col77[9]),
        .b(stage2_col77[10]),
        .c_in(stage2_col77[11]),
        .s(fa_s2_c77_n207_s),
        .c_out(fa_s2_c77_n207_c)
    );

    fa fa_s2_c77_n208 (
        .a(stage2_col77[12]),
        .b(stage2_col77[13]),
        .c_in(stage2_col77[14]),
        .s(fa_s2_c77_n208_s),
        .c_out(fa_s2_c77_n208_c)
    );

    fa fa_s2_c78_n209 (
        .a(stage2_col78[0]),
        .b(stage2_col78[1]),
        .c_in(stage2_col78[2]),
        .s(fa_s2_c78_n209_s),
        .c_out(fa_s2_c78_n209_c)
    );

    fa fa_s2_c78_n210 (
        .a(stage2_col78[3]),
        .b(stage2_col78[4]),
        .c_in(stage2_col78[5]),
        .s(fa_s2_c78_n210_s),
        .c_out(fa_s2_c78_n210_c)
    );

    fa fa_s2_c78_n211 (
        .a(stage2_col78[6]),
        .b(stage2_col78[7]),
        .c_in(stage2_col78[8]),
        .s(fa_s2_c78_n211_s),
        .c_out(fa_s2_c78_n211_c)
    );

    fa fa_s2_c78_n212 (
        .a(stage2_col78[9]),
        .b(stage2_col78[10]),
        .c_in(stage2_col78[11]),
        .s(fa_s2_c78_n212_s),
        .c_out(fa_s2_c78_n212_c)
    );

    fa fa_s2_c79_n213 (
        .a(stage2_col79[0]),
        .b(stage2_col79[1]),
        .c_in(stage2_col79[2]),
        .s(fa_s2_c79_n213_s),
        .c_out(fa_s2_c79_n213_c)
    );

    fa fa_s2_c79_n214 (
        .a(stage2_col79[3]),
        .b(stage2_col79[4]),
        .c_in(stage2_col79[5]),
        .s(fa_s2_c79_n214_s),
        .c_out(fa_s2_c79_n214_c)
    );

    fa fa_s2_c79_n215 (
        .a(stage2_col79[6]),
        .b(stage2_col79[7]),
        .c_in(stage2_col79[8]),
        .s(fa_s2_c79_n215_s),
        .c_out(fa_s2_c79_n215_c)
    );

    fa fa_s2_c79_n216 (
        .a(stage2_col79[9]),
        .b(stage2_col79[10]),
        .c_in(stage2_col79[11]),
        .s(fa_s2_c79_n216_s),
        .c_out(fa_s2_c79_n216_c)
    );

    fa fa_s2_c79_n217 (
        .a(stage2_col79[12]),
        .b(stage2_col79[13]),
        .c_in(stage2_col79[14]),
        .s(fa_s2_c79_n217_s),
        .c_out(fa_s2_c79_n217_c)
    );

    fa fa_s2_c80_n218 (
        .a(stage2_col80[0]),
        .b(stage2_col80[1]),
        .c_in(stage2_col80[2]),
        .s(fa_s2_c80_n218_s),
        .c_out(fa_s2_c80_n218_c)
    );

    fa fa_s2_c80_n219 (
        .a(stage2_col80[3]),
        .b(stage2_col80[4]),
        .c_in(stage2_col80[5]),
        .s(fa_s2_c80_n219_s),
        .c_out(fa_s2_c80_n219_c)
    );

    fa fa_s2_c80_n220 (
        .a(stage2_col80[6]),
        .b(stage2_col80[7]),
        .c_in(stage2_col80[8]),
        .s(fa_s2_c80_n220_s),
        .c_out(fa_s2_c80_n220_c)
    );

    fa fa_s2_c80_n221 (
        .a(stage2_col80[9]),
        .b(stage2_col80[10]),
        .c_in(stage2_col80[11]),
        .s(fa_s2_c80_n221_s),
        .c_out(fa_s2_c80_n221_c)
    );

    fa fa_s2_c81_n222 (
        .a(stage2_col81[0]),
        .b(stage2_col81[1]),
        .c_in(stage2_col81[2]),
        .s(fa_s2_c81_n222_s),
        .c_out(fa_s2_c81_n222_c)
    );

    fa fa_s2_c81_n223 (
        .a(stage2_col81[3]),
        .b(stage2_col81[4]),
        .c_in(stage2_col81[5]),
        .s(fa_s2_c81_n223_s),
        .c_out(fa_s2_c81_n223_c)
    );

    fa fa_s2_c81_n224 (
        .a(stage2_col81[6]),
        .b(stage2_col81[7]),
        .c_in(stage2_col81[8]),
        .s(fa_s2_c81_n224_s),
        .c_out(fa_s2_c81_n224_c)
    );

    fa fa_s2_c81_n225 (
        .a(stage2_col81[9]),
        .b(stage2_col81[10]),
        .c_in(stage2_col81[11]),
        .s(fa_s2_c81_n225_s),
        .c_out(fa_s2_c81_n225_c)
    );

    fa fa_s2_c81_n226 (
        .a(stage2_col81[12]),
        .b(stage2_col81[13]),
        .c_in(stage2_col81[14]),
        .s(fa_s2_c81_n226_s),
        .c_out(fa_s2_c81_n226_c)
    );

    fa fa_s2_c82_n227 (
        .a(stage2_col82[0]),
        .b(stage2_col82[1]),
        .c_in(stage2_col82[2]),
        .s(fa_s2_c82_n227_s),
        .c_out(fa_s2_c82_n227_c)
    );

    fa fa_s2_c82_n228 (
        .a(stage2_col82[3]),
        .b(stage2_col82[4]),
        .c_in(stage2_col82[5]),
        .s(fa_s2_c82_n228_s),
        .c_out(fa_s2_c82_n228_c)
    );

    fa fa_s2_c82_n229 (
        .a(stage2_col82[6]),
        .b(stage2_col82[7]),
        .c_in(stage2_col82[8]),
        .s(fa_s2_c82_n229_s),
        .c_out(fa_s2_c82_n229_c)
    );

    fa fa_s2_c82_n230 (
        .a(stage2_col82[9]),
        .b(stage2_col82[10]),
        .c_in(stage2_col82[11]),
        .s(fa_s2_c82_n230_s),
        .c_out(fa_s2_c82_n230_c)
    );

    fa fa_s2_c83_n231 (
        .a(stage2_col83[0]),
        .b(stage2_col83[1]),
        .c_in(stage2_col83[2]),
        .s(fa_s2_c83_n231_s),
        .c_out(fa_s2_c83_n231_c)
    );

    fa fa_s2_c83_n232 (
        .a(stage2_col83[3]),
        .b(stage2_col83[4]),
        .c_in(stage2_col83[5]),
        .s(fa_s2_c83_n232_s),
        .c_out(fa_s2_c83_n232_c)
    );

    fa fa_s2_c83_n233 (
        .a(stage2_col83[6]),
        .b(stage2_col83[7]),
        .c_in(stage2_col83[8]),
        .s(fa_s2_c83_n233_s),
        .c_out(fa_s2_c83_n233_c)
    );

    fa fa_s2_c83_n234 (
        .a(stage2_col83[9]),
        .b(stage2_col83[10]),
        .c_in(stage2_col83[11]),
        .s(fa_s2_c83_n234_s),
        .c_out(fa_s2_c83_n234_c)
    );

    fa fa_s2_c83_n235 (
        .a(stage2_col83[12]),
        .b(stage2_col83[13]),
        .c_in(stage2_col83[14]),
        .s(fa_s2_c83_n235_s),
        .c_out(fa_s2_c83_n235_c)
    );

    fa fa_s2_c84_n236 (
        .a(stage2_col84[0]),
        .b(stage2_col84[1]),
        .c_in(stage2_col84[2]),
        .s(fa_s2_c84_n236_s),
        .c_out(fa_s2_c84_n236_c)
    );

    fa fa_s2_c84_n237 (
        .a(stage2_col84[3]),
        .b(stage2_col84[4]),
        .c_in(stage2_col84[5]),
        .s(fa_s2_c84_n237_s),
        .c_out(fa_s2_c84_n237_c)
    );

    fa fa_s2_c84_n238 (
        .a(stage2_col84[6]),
        .b(stage2_col84[7]),
        .c_in(stage2_col84[8]),
        .s(fa_s2_c84_n238_s),
        .c_out(fa_s2_c84_n238_c)
    );

    fa fa_s2_c84_n239 (
        .a(stage2_col84[9]),
        .b(stage2_col84[10]),
        .c_in(stage2_col84[11]),
        .s(fa_s2_c84_n239_s),
        .c_out(fa_s2_c84_n239_c)
    );

    fa fa_s2_c85_n240 (
        .a(stage2_col85[0]),
        .b(stage2_col85[1]),
        .c_in(stage2_col85[2]),
        .s(fa_s2_c85_n240_s),
        .c_out(fa_s2_c85_n240_c)
    );

    fa fa_s2_c85_n241 (
        .a(stage2_col85[3]),
        .b(stage2_col85[4]),
        .c_in(stage2_col85[5]),
        .s(fa_s2_c85_n241_s),
        .c_out(fa_s2_c85_n241_c)
    );

    fa fa_s2_c85_n242 (
        .a(stage2_col85[6]),
        .b(stage2_col85[7]),
        .c_in(stage2_col85[8]),
        .s(fa_s2_c85_n242_s),
        .c_out(fa_s2_c85_n242_c)
    );

    fa fa_s2_c85_n243 (
        .a(stage2_col85[9]),
        .b(stage2_col85[10]),
        .c_in(stage2_col85[11]),
        .s(fa_s2_c85_n243_s),
        .c_out(fa_s2_c85_n243_c)
    );

    fa fa_s2_c85_n244 (
        .a(stage2_col85[12]),
        .b(stage2_col85[13]),
        .c_in(stage2_col85[14]),
        .s(fa_s2_c85_n244_s),
        .c_out(fa_s2_c85_n244_c)
    );

    fa fa_s2_c86_n245 (
        .a(stage2_col86[0]),
        .b(stage2_col86[1]),
        .c_in(stage2_col86[2]),
        .s(fa_s2_c86_n245_s),
        .c_out(fa_s2_c86_n245_c)
    );

    fa fa_s2_c86_n246 (
        .a(stage2_col86[3]),
        .b(stage2_col86[4]),
        .c_in(stage2_col86[5]),
        .s(fa_s2_c86_n246_s),
        .c_out(fa_s2_c86_n246_c)
    );

    fa fa_s2_c86_n247 (
        .a(stage2_col86[6]),
        .b(stage2_col86[7]),
        .c_in(stage2_col86[8]),
        .s(fa_s2_c86_n247_s),
        .c_out(fa_s2_c86_n247_c)
    );

    fa fa_s2_c86_n248 (
        .a(stage2_col86[9]),
        .b(stage2_col86[10]),
        .c_in(stage2_col86[11]),
        .s(fa_s2_c86_n248_s),
        .c_out(fa_s2_c86_n248_c)
    );

    fa fa_s2_c87_n249 (
        .a(stage2_col87[0]),
        .b(stage2_col87[1]),
        .c_in(stage2_col87[2]),
        .s(fa_s2_c87_n249_s),
        .c_out(fa_s2_c87_n249_c)
    );

    fa fa_s2_c87_n250 (
        .a(stage2_col87[3]),
        .b(stage2_col87[4]),
        .c_in(stage2_col87[5]),
        .s(fa_s2_c87_n250_s),
        .c_out(fa_s2_c87_n250_c)
    );

    fa fa_s2_c87_n251 (
        .a(stage2_col87[6]),
        .b(stage2_col87[7]),
        .c_in(stage2_col87[8]),
        .s(fa_s2_c87_n251_s),
        .c_out(fa_s2_c87_n251_c)
    );

    fa fa_s2_c87_n252 (
        .a(stage2_col87[9]),
        .b(stage2_col87[10]),
        .c_in(stage2_col87[11]),
        .s(fa_s2_c87_n252_s),
        .c_out(fa_s2_c87_n252_c)
    );

    fa fa_s2_c87_n253 (
        .a(stage2_col87[12]),
        .b(stage2_col87[13]),
        .c_in(stage2_col87[14]),
        .s(fa_s2_c87_n253_s),
        .c_out(fa_s2_c87_n253_c)
    );

    fa fa_s2_c88_n254 (
        .a(stage2_col88[0]),
        .b(stage2_col88[1]),
        .c_in(stage2_col88[2]),
        .s(fa_s2_c88_n254_s),
        .c_out(fa_s2_c88_n254_c)
    );

    fa fa_s2_c88_n255 (
        .a(stage2_col88[3]),
        .b(stage2_col88[4]),
        .c_in(stage2_col88[5]),
        .s(fa_s2_c88_n255_s),
        .c_out(fa_s2_c88_n255_c)
    );

    fa fa_s2_c88_n256 (
        .a(stage2_col88[6]),
        .b(stage2_col88[7]),
        .c_in(stage2_col88[8]),
        .s(fa_s2_c88_n256_s),
        .c_out(fa_s2_c88_n256_c)
    );

    fa fa_s2_c88_n257 (
        .a(stage2_col88[9]),
        .b(stage2_col88[10]),
        .c_in(stage2_col88[11]),
        .s(fa_s2_c88_n257_s),
        .c_out(fa_s2_c88_n257_c)
    );

    fa fa_s2_c89_n258 (
        .a(stage2_col89[0]),
        .b(stage2_col89[1]),
        .c_in(stage2_col89[2]),
        .s(fa_s2_c89_n258_s),
        .c_out(fa_s2_c89_n258_c)
    );

    fa fa_s2_c89_n259 (
        .a(stage2_col89[3]),
        .b(stage2_col89[4]),
        .c_in(stage2_col89[5]),
        .s(fa_s2_c89_n259_s),
        .c_out(fa_s2_c89_n259_c)
    );

    fa fa_s2_c89_n260 (
        .a(stage2_col89[6]),
        .b(stage2_col89[7]),
        .c_in(stage2_col89[8]),
        .s(fa_s2_c89_n260_s),
        .c_out(fa_s2_c89_n260_c)
    );

    fa fa_s2_c89_n261 (
        .a(stage2_col89[9]),
        .b(stage2_col89[10]),
        .c_in(stage2_col89[11]),
        .s(fa_s2_c89_n261_s),
        .c_out(fa_s2_c89_n261_c)
    );

    fa fa_s2_c89_n262 (
        .a(stage2_col89[12]),
        .b(stage2_col89[13]),
        .c_in(stage2_col89[14]),
        .s(fa_s2_c89_n262_s),
        .c_out(fa_s2_c89_n262_c)
    );

    fa fa_s2_c90_n263 (
        .a(stage2_col90[0]),
        .b(stage2_col90[1]),
        .c_in(stage2_col90[2]),
        .s(fa_s2_c90_n263_s),
        .c_out(fa_s2_c90_n263_c)
    );

    fa fa_s2_c90_n264 (
        .a(stage2_col90[3]),
        .b(stage2_col90[4]),
        .c_in(stage2_col90[5]),
        .s(fa_s2_c90_n264_s),
        .c_out(fa_s2_c90_n264_c)
    );

    fa fa_s2_c90_n265 (
        .a(stage2_col90[6]),
        .b(stage2_col90[7]),
        .c_in(stage2_col90[8]),
        .s(fa_s2_c90_n265_s),
        .c_out(fa_s2_c90_n265_c)
    );

    fa fa_s2_c90_n266 (
        .a(stage2_col90[9]),
        .b(stage2_col90[10]),
        .c_in(stage2_col90[11]),
        .s(fa_s2_c90_n266_s),
        .c_out(fa_s2_c90_n266_c)
    );

    fa fa_s2_c91_n267 (
        .a(stage2_col91[0]),
        .b(stage2_col91[1]),
        .c_in(stage2_col91[2]),
        .s(fa_s2_c91_n267_s),
        .c_out(fa_s2_c91_n267_c)
    );

    fa fa_s2_c91_n268 (
        .a(stage2_col91[3]),
        .b(stage2_col91[4]),
        .c_in(stage2_col91[5]),
        .s(fa_s2_c91_n268_s),
        .c_out(fa_s2_c91_n268_c)
    );

    fa fa_s2_c91_n269 (
        .a(stage2_col91[6]),
        .b(stage2_col91[7]),
        .c_in(stage2_col91[8]),
        .s(fa_s2_c91_n269_s),
        .c_out(fa_s2_c91_n269_c)
    );

    fa fa_s2_c91_n270 (
        .a(stage2_col91[9]),
        .b(stage2_col91[10]),
        .c_in(stage2_col91[11]),
        .s(fa_s2_c91_n270_s),
        .c_out(fa_s2_c91_n270_c)
    );

    fa fa_s2_c91_n271 (
        .a(stage2_col91[12]),
        .b(stage2_col91[13]),
        .c_in(stage2_col91[14]),
        .s(fa_s2_c91_n271_s),
        .c_out(fa_s2_c91_n271_c)
    );

    fa fa_s2_c92_n272 (
        .a(stage2_col92[0]),
        .b(stage2_col92[1]),
        .c_in(stage2_col92[2]),
        .s(fa_s2_c92_n272_s),
        .c_out(fa_s2_c92_n272_c)
    );

    fa fa_s2_c92_n273 (
        .a(stage2_col92[3]),
        .b(stage2_col92[4]),
        .c_in(stage2_col92[5]),
        .s(fa_s2_c92_n273_s),
        .c_out(fa_s2_c92_n273_c)
    );

    fa fa_s2_c92_n274 (
        .a(stage2_col92[6]),
        .b(stage2_col92[7]),
        .c_in(stage2_col92[8]),
        .s(fa_s2_c92_n274_s),
        .c_out(fa_s2_c92_n274_c)
    );

    fa fa_s2_c92_n275 (
        .a(stage2_col92[9]),
        .b(stage2_col92[10]),
        .c_in(stage2_col92[11]),
        .s(fa_s2_c92_n275_s),
        .c_out(fa_s2_c92_n275_c)
    );

    fa fa_s2_c93_n276 (
        .a(stage2_col93[0]),
        .b(stage2_col93[1]),
        .c_in(stage2_col93[2]),
        .s(fa_s2_c93_n276_s),
        .c_out(fa_s2_c93_n276_c)
    );

    fa fa_s2_c93_n277 (
        .a(stage2_col93[3]),
        .b(stage2_col93[4]),
        .c_in(stage2_col93[5]),
        .s(fa_s2_c93_n277_s),
        .c_out(fa_s2_c93_n277_c)
    );

    fa fa_s2_c93_n278 (
        .a(stage2_col93[6]),
        .b(stage2_col93[7]),
        .c_in(stage2_col93[8]),
        .s(fa_s2_c93_n278_s),
        .c_out(fa_s2_c93_n278_c)
    );

    fa fa_s2_c93_n279 (
        .a(stage2_col93[9]),
        .b(stage2_col93[10]),
        .c_in(stage2_col93[11]),
        .s(fa_s2_c93_n279_s),
        .c_out(fa_s2_c93_n279_c)
    );

    fa fa_s2_c93_n280 (
        .a(stage2_col93[12]),
        .b(stage2_col93[13]),
        .c_in(stage2_col93[14]),
        .s(fa_s2_c93_n280_s),
        .c_out(fa_s2_c93_n280_c)
    );

    fa fa_s2_c94_n281 (
        .a(stage2_col94[0]),
        .b(stage2_col94[1]),
        .c_in(stage2_col94[2]),
        .s(fa_s2_c94_n281_s),
        .c_out(fa_s2_c94_n281_c)
    );

    fa fa_s2_c94_n282 (
        .a(stage2_col94[3]),
        .b(stage2_col94[4]),
        .c_in(stage2_col94[5]),
        .s(fa_s2_c94_n282_s),
        .c_out(fa_s2_c94_n282_c)
    );

    fa fa_s2_c94_n283 (
        .a(stage2_col94[6]),
        .b(stage2_col94[7]),
        .c_in(stage2_col94[8]),
        .s(fa_s2_c94_n283_s),
        .c_out(fa_s2_c94_n283_c)
    );

    fa fa_s2_c94_n284 (
        .a(stage2_col94[9]),
        .b(stage2_col94[10]),
        .c_in(stage2_col94[11]),
        .s(fa_s2_c94_n284_s),
        .c_out(fa_s2_c94_n284_c)
    );

    fa fa_s2_c95_n285 (
        .a(stage2_col95[0]),
        .b(stage2_col95[1]),
        .c_in(stage2_col95[2]),
        .s(fa_s2_c95_n285_s),
        .c_out(fa_s2_c95_n285_c)
    );

    fa fa_s2_c95_n286 (
        .a(stage2_col95[3]),
        .b(stage2_col95[4]),
        .c_in(stage2_col95[5]),
        .s(fa_s2_c95_n286_s),
        .c_out(fa_s2_c95_n286_c)
    );

    fa fa_s2_c95_n287 (
        .a(stage2_col95[6]),
        .b(stage2_col95[7]),
        .c_in(stage2_col95[8]),
        .s(fa_s2_c95_n287_s),
        .c_out(fa_s2_c95_n287_c)
    );

    fa fa_s2_c95_n288 (
        .a(stage2_col95[9]),
        .b(stage2_col95[10]),
        .c_in(stage2_col95[11]),
        .s(fa_s2_c95_n288_s),
        .c_out(fa_s2_c95_n288_c)
    );

    fa fa_s2_c95_n289 (
        .a(stage2_col95[12]),
        .b(stage2_col95[13]),
        .c_in(stage2_col95[14]),
        .s(fa_s2_c95_n289_s),
        .c_out(fa_s2_c95_n289_c)
    );

    fa fa_s2_c96_n290 (
        .a(stage2_col96[0]),
        .b(stage2_col96[1]),
        .c_in(stage2_col96[2]),
        .s(fa_s2_c96_n290_s),
        .c_out(fa_s2_c96_n290_c)
    );

    fa fa_s2_c96_n291 (
        .a(stage2_col96[3]),
        .b(stage2_col96[4]),
        .c_in(stage2_col96[5]),
        .s(fa_s2_c96_n291_s),
        .c_out(fa_s2_c96_n291_c)
    );

    fa fa_s2_c96_n292 (
        .a(stage2_col96[6]),
        .b(stage2_col96[7]),
        .c_in(stage2_col96[8]),
        .s(fa_s2_c96_n292_s),
        .c_out(fa_s2_c96_n292_c)
    );

    fa fa_s2_c96_n293 (
        .a(stage2_col96[9]),
        .b(stage2_col96[10]),
        .c_in(stage2_col96[11]),
        .s(fa_s2_c96_n293_s),
        .c_out(fa_s2_c96_n293_c)
    );

    fa fa_s2_c97_n294 (
        .a(stage2_col97[0]),
        .b(stage2_col97[1]),
        .c_in(stage2_col97[2]),
        .s(fa_s2_c97_n294_s),
        .c_out(fa_s2_c97_n294_c)
    );

    fa fa_s2_c97_n295 (
        .a(stage2_col97[3]),
        .b(stage2_col97[4]),
        .c_in(stage2_col97[5]),
        .s(fa_s2_c97_n295_s),
        .c_out(fa_s2_c97_n295_c)
    );

    fa fa_s2_c97_n296 (
        .a(stage2_col97[6]),
        .b(stage2_col97[7]),
        .c_in(stage2_col97[8]),
        .s(fa_s2_c97_n296_s),
        .c_out(fa_s2_c97_n296_c)
    );

    fa fa_s2_c97_n297 (
        .a(stage2_col97[9]),
        .b(stage2_col97[10]),
        .c_in(stage2_col97[11]),
        .s(fa_s2_c97_n297_s),
        .c_out(fa_s2_c97_n297_c)
    );

    fa fa_s2_c97_n298 (
        .a(stage2_col97[12]),
        .b(stage2_col97[13]),
        .c_in(stage2_col97[14]),
        .s(fa_s2_c97_n298_s),
        .c_out(fa_s2_c97_n298_c)
    );

    fa fa_s2_c98_n299 (
        .a(stage2_col98[0]),
        .b(stage2_col98[1]),
        .c_in(stage2_col98[2]),
        .s(fa_s2_c98_n299_s),
        .c_out(fa_s2_c98_n299_c)
    );

    fa fa_s2_c98_n300 (
        .a(stage2_col98[3]),
        .b(stage2_col98[4]),
        .c_in(stage2_col98[5]),
        .s(fa_s2_c98_n300_s),
        .c_out(fa_s2_c98_n300_c)
    );

    fa fa_s2_c98_n301 (
        .a(stage2_col98[6]),
        .b(stage2_col98[7]),
        .c_in(stage2_col98[8]),
        .s(fa_s2_c98_n301_s),
        .c_out(fa_s2_c98_n301_c)
    );

    fa fa_s2_c98_n302 (
        .a(stage2_col98[9]),
        .b(stage2_col98[10]),
        .c_in(stage2_col98[11]),
        .s(fa_s2_c98_n302_s),
        .c_out(fa_s2_c98_n302_c)
    );

    fa fa_s2_c99_n303 (
        .a(stage2_col99[0]),
        .b(stage2_col99[1]),
        .c_in(stage2_col99[2]),
        .s(fa_s2_c99_n303_s),
        .c_out(fa_s2_c99_n303_c)
    );

    fa fa_s2_c99_n304 (
        .a(stage2_col99[3]),
        .b(stage2_col99[4]),
        .c_in(stage2_col99[5]),
        .s(fa_s2_c99_n304_s),
        .c_out(fa_s2_c99_n304_c)
    );

    fa fa_s2_c99_n305 (
        .a(stage2_col99[6]),
        .b(stage2_col99[7]),
        .c_in(stage2_col99[8]),
        .s(fa_s2_c99_n305_s),
        .c_out(fa_s2_c99_n305_c)
    );

    fa fa_s2_c99_n306 (
        .a(stage2_col99[9]),
        .b(stage2_col99[10]),
        .c_in(stage2_col99[11]),
        .s(fa_s2_c99_n306_s),
        .c_out(fa_s2_c99_n306_c)
    );

    fa fa_s2_c99_n307 (
        .a(stage2_col99[12]),
        .b(stage2_col99[13]),
        .c_in(stage2_col99[14]),
        .s(fa_s2_c99_n307_s),
        .c_out(fa_s2_c99_n307_c)
    );

    fa fa_s2_c100_n308 (
        .a(stage2_col100[0]),
        .b(stage2_col100[1]),
        .c_in(stage2_col100[2]),
        .s(fa_s2_c100_n308_s),
        .c_out(fa_s2_c100_n308_c)
    );

    fa fa_s2_c100_n309 (
        .a(stage2_col100[3]),
        .b(stage2_col100[4]),
        .c_in(stage2_col100[5]),
        .s(fa_s2_c100_n309_s),
        .c_out(fa_s2_c100_n309_c)
    );

    fa fa_s2_c100_n310 (
        .a(stage2_col100[6]),
        .b(stage2_col100[7]),
        .c_in(stage2_col100[8]),
        .s(fa_s2_c100_n310_s),
        .c_out(fa_s2_c100_n310_c)
    );

    fa fa_s2_c100_n311 (
        .a(stage2_col100[9]),
        .b(stage2_col100[10]),
        .c_in(stage2_col100[11]),
        .s(fa_s2_c100_n311_s),
        .c_out(fa_s2_c100_n311_c)
    );

    fa fa_s2_c101_n312 (
        .a(stage2_col101[0]),
        .b(stage2_col101[1]),
        .c_in(stage2_col101[2]),
        .s(fa_s2_c101_n312_s),
        .c_out(fa_s2_c101_n312_c)
    );

    fa fa_s2_c101_n313 (
        .a(stage2_col101[3]),
        .b(stage2_col101[4]),
        .c_in(stage2_col101[5]),
        .s(fa_s2_c101_n313_s),
        .c_out(fa_s2_c101_n313_c)
    );

    fa fa_s2_c101_n314 (
        .a(stage2_col101[6]),
        .b(stage2_col101[7]),
        .c_in(stage2_col101[8]),
        .s(fa_s2_c101_n314_s),
        .c_out(fa_s2_c101_n314_c)
    );

    fa fa_s2_c101_n315 (
        .a(stage2_col101[9]),
        .b(stage2_col101[10]),
        .c_in(stage2_col101[11]),
        .s(fa_s2_c101_n315_s),
        .c_out(fa_s2_c101_n315_c)
    );

    fa fa_s2_c101_n316 (
        .a(stage2_col101[12]),
        .b(stage2_col101[13]),
        .c_in(stage2_col101[14]),
        .s(fa_s2_c101_n316_s),
        .c_out(fa_s2_c101_n316_c)
    );

    fa fa_s2_c102_n317 (
        .a(stage2_col102[0]),
        .b(stage2_col102[1]),
        .c_in(stage2_col102[2]),
        .s(fa_s2_c102_n317_s),
        .c_out(fa_s2_c102_n317_c)
    );

    fa fa_s2_c102_n318 (
        .a(stage2_col102[3]),
        .b(stage2_col102[4]),
        .c_in(stage2_col102[5]),
        .s(fa_s2_c102_n318_s),
        .c_out(fa_s2_c102_n318_c)
    );

    fa fa_s2_c102_n319 (
        .a(stage2_col102[6]),
        .b(stage2_col102[7]),
        .c_in(stage2_col102[8]),
        .s(fa_s2_c102_n319_s),
        .c_out(fa_s2_c102_n319_c)
    );

    fa fa_s2_c102_n320 (
        .a(stage2_col102[9]),
        .b(stage2_col102[10]),
        .c_in(stage2_col102[11]),
        .s(fa_s2_c102_n320_s),
        .c_out(fa_s2_c102_n320_c)
    );

    fa fa_s2_c103_n321 (
        .a(stage2_col103[0]),
        .b(stage2_col103[1]),
        .c_in(stage2_col103[2]),
        .s(fa_s2_c103_n321_s),
        .c_out(fa_s2_c103_n321_c)
    );

    fa fa_s2_c103_n322 (
        .a(stage2_col103[3]),
        .b(stage2_col103[4]),
        .c_in(stage2_col103[5]),
        .s(fa_s2_c103_n322_s),
        .c_out(fa_s2_c103_n322_c)
    );

    fa fa_s2_c103_n323 (
        .a(stage2_col103[6]),
        .b(stage2_col103[7]),
        .c_in(stage2_col103[8]),
        .s(fa_s2_c103_n323_s),
        .c_out(fa_s2_c103_n323_c)
    );

    fa fa_s2_c103_n324 (
        .a(stage2_col103[9]),
        .b(stage2_col103[10]),
        .c_in(stage2_col103[11]),
        .s(fa_s2_c103_n324_s),
        .c_out(fa_s2_c103_n324_c)
    );

    fa fa_s2_c103_n325 (
        .a(stage2_col103[12]),
        .b(stage2_col103[13]),
        .c_in(stage2_col103[14]),
        .s(fa_s2_c103_n325_s),
        .c_out(fa_s2_c103_n325_c)
    );

    fa fa_s2_c104_n326 (
        .a(stage2_col104[0]),
        .b(stage2_col104[1]),
        .c_in(stage2_col104[2]),
        .s(fa_s2_c104_n326_s),
        .c_out(fa_s2_c104_n326_c)
    );

    fa fa_s2_c104_n327 (
        .a(stage2_col104[3]),
        .b(stage2_col104[4]),
        .c_in(stage2_col104[5]),
        .s(fa_s2_c104_n327_s),
        .c_out(fa_s2_c104_n327_c)
    );

    fa fa_s2_c104_n328 (
        .a(stage2_col104[6]),
        .b(stage2_col104[7]),
        .c_in(stage2_col104[8]),
        .s(fa_s2_c104_n328_s),
        .c_out(fa_s2_c104_n328_c)
    );

    fa fa_s2_c104_n329 (
        .a(stage2_col104[9]),
        .b(stage2_col104[10]),
        .c_in(stage2_col104[11]),
        .s(fa_s2_c104_n329_s),
        .c_out(fa_s2_c104_n329_c)
    );

    fa fa_s2_c105_n330 (
        .a(stage2_col105[0]),
        .b(stage2_col105[1]),
        .c_in(stage2_col105[2]),
        .s(fa_s2_c105_n330_s),
        .c_out(fa_s2_c105_n330_c)
    );

    fa fa_s2_c105_n331 (
        .a(stage2_col105[3]),
        .b(stage2_col105[4]),
        .c_in(stage2_col105[5]),
        .s(fa_s2_c105_n331_s),
        .c_out(fa_s2_c105_n331_c)
    );

    fa fa_s2_c105_n332 (
        .a(stage2_col105[6]),
        .b(stage2_col105[7]),
        .c_in(stage2_col105[8]),
        .s(fa_s2_c105_n332_s),
        .c_out(fa_s2_c105_n332_c)
    );

    fa fa_s2_c105_n333 (
        .a(stage2_col105[9]),
        .b(stage2_col105[10]),
        .c_in(stage2_col105[11]),
        .s(fa_s2_c105_n333_s),
        .c_out(fa_s2_c105_n333_c)
    );

    fa fa_s2_c105_n334 (
        .a(stage2_col105[12]),
        .b(stage2_col105[13]),
        .c_in(stage2_col105[14]),
        .s(fa_s2_c105_n334_s),
        .c_out(fa_s2_c105_n334_c)
    );

    fa fa_s2_c106_n335 (
        .a(stage2_col106[0]),
        .b(stage2_col106[1]),
        .c_in(stage2_col106[2]),
        .s(fa_s2_c106_n335_s),
        .c_out(fa_s2_c106_n335_c)
    );

    fa fa_s2_c106_n336 (
        .a(stage2_col106[3]),
        .b(stage2_col106[4]),
        .c_in(stage2_col106[5]),
        .s(fa_s2_c106_n336_s),
        .c_out(fa_s2_c106_n336_c)
    );

    fa fa_s2_c106_n337 (
        .a(stage2_col106[6]),
        .b(stage2_col106[7]),
        .c_in(stage2_col106[8]),
        .s(fa_s2_c106_n337_s),
        .c_out(fa_s2_c106_n337_c)
    );

    fa fa_s2_c106_n338 (
        .a(stage2_col106[9]),
        .b(stage2_col106[10]),
        .c_in(stage2_col106[11]),
        .s(fa_s2_c106_n338_s),
        .c_out(fa_s2_c106_n338_c)
    );

    fa fa_s2_c107_n339 (
        .a(stage2_col107[0]),
        .b(stage2_col107[1]),
        .c_in(stage2_col107[2]),
        .s(fa_s2_c107_n339_s),
        .c_out(fa_s2_c107_n339_c)
    );

    fa fa_s2_c107_n340 (
        .a(stage2_col107[3]),
        .b(stage2_col107[4]),
        .c_in(stage2_col107[5]),
        .s(fa_s2_c107_n340_s),
        .c_out(fa_s2_c107_n340_c)
    );

    fa fa_s2_c107_n341 (
        .a(stage2_col107[6]),
        .b(stage2_col107[7]),
        .c_in(stage2_col107[8]),
        .s(fa_s2_c107_n341_s),
        .c_out(fa_s2_c107_n341_c)
    );

    fa fa_s2_c107_n342 (
        .a(stage2_col107[9]),
        .b(stage2_col107[10]),
        .c_in(stage2_col107[11]),
        .s(fa_s2_c107_n342_s),
        .c_out(fa_s2_c107_n342_c)
    );

    fa fa_s2_c107_n343 (
        .a(stage2_col107[12]),
        .b(stage2_col107[13]),
        .c_in(stage2_col107[14]),
        .s(fa_s2_c107_n343_s),
        .c_out(fa_s2_c107_n343_c)
    );

    fa fa_s2_c108_n344 (
        .a(stage2_col108[0]),
        .b(stage2_col108[1]),
        .c_in(stage2_col108[2]),
        .s(fa_s2_c108_n344_s),
        .c_out(fa_s2_c108_n344_c)
    );

    fa fa_s2_c108_n345 (
        .a(stage2_col108[3]),
        .b(stage2_col108[4]),
        .c_in(stage2_col108[5]),
        .s(fa_s2_c108_n345_s),
        .c_out(fa_s2_c108_n345_c)
    );

    fa fa_s2_c108_n346 (
        .a(stage2_col108[6]),
        .b(stage2_col108[7]),
        .c_in(stage2_col108[8]),
        .s(fa_s2_c108_n346_s),
        .c_out(fa_s2_c108_n346_c)
    );

    fa fa_s2_c108_n347 (
        .a(stage2_col108[9]),
        .b(stage2_col108[10]),
        .c_in(stage2_col108[11]),
        .s(fa_s2_c108_n347_s),
        .c_out(fa_s2_c108_n347_c)
    );

    fa fa_s2_c109_n348 (
        .a(stage2_col109[0]),
        .b(stage2_col109[1]),
        .c_in(stage2_col109[2]),
        .s(fa_s2_c109_n348_s),
        .c_out(fa_s2_c109_n348_c)
    );

    fa fa_s2_c109_n349 (
        .a(stage2_col109[3]),
        .b(stage2_col109[4]),
        .c_in(stage2_col109[5]),
        .s(fa_s2_c109_n349_s),
        .c_out(fa_s2_c109_n349_c)
    );

    fa fa_s2_c109_n350 (
        .a(stage2_col109[6]),
        .b(stage2_col109[7]),
        .c_in(stage2_col109[8]),
        .s(fa_s2_c109_n350_s),
        .c_out(fa_s2_c109_n350_c)
    );

    fa fa_s2_c109_n351 (
        .a(stage2_col109[9]),
        .b(stage2_col109[10]),
        .c_in(stage2_col109[11]),
        .s(fa_s2_c109_n351_s),
        .c_out(fa_s2_c109_n351_c)
    );

    fa fa_s2_c109_n352 (
        .a(stage2_col109[12]),
        .b(stage2_col109[13]),
        .c_in(stage2_col109[14]),
        .s(fa_s2_c109_n352_s),
        .c_out(fa_s2_c109_n352_c)
    );

    fa fa_s2_c110_n353 (
        .a(stage2_col110[0]),
        .b(stage2_col110[1]),
        .c_in(stage2_col110[2]),
        .s(fa_s2_c110_n353_s),
        .c_out(fa_s2_c110_n353_c)
    );

    fa fa_s2_c110_n354 (
        .a(stage2_col110[3]),
        .b(stage2_col110[4]),
        .c_in(stage2_col110[5]),
        .s(fa_s2_c110_n354_s),
        .c_out(fa_s2_c110_n354_c)
    );

    fa fa_s2_c110_n355 (
        .a(stage2_col110[6]),
        .b(stage2_col110[7]),
        .c_in(stage2_col110[8]),
        .s(fa_s2_c110_n355_s),
        .c_out(fa_s2_c110_n355_c)
    );

    fa fa_s2_c110_n356 (
        .a(stage2_col110[9]),
        .b(stage2_col110[10]),
        .c_in(stage2_col110[11]),
        .s(fa_s2_c110_n356_s),
        .c_out(fa_s2_c110_n356_c)
    );

    fa fa_s2_c111_n357 (
        .a(stage2_col111[0]),
        .b(stage2_col111[1]),
        .c_in(stage2_col111[2]),
        .s(fa_s2_c111_n357_s),
        .c_out(fa_s2_c111_n357_c)
    );

    fa fa_s2_c111_n358 (
        .a(stage2_col111[3]),
        .b(stage2_col111[4]),
        .c_in(stage2_col111[5]),
        .s(fa_s2_c111_n358_s),
        .c_out(fa_s2_c111_n358_c)
    );

    fa fa_s2_c111_n359 (
        .a(stage2_col111[6]),
        .b(stage2_col111[7]),
        .c_in(stage2_col111[8]),
        .s(fa_s2_c111_n359_s),
        .c_out(fa_s2_c111_n359_c)
    );

    fa fa_s2_c111_n360 (
        .a(stage2_col111[9]),
        .b(stage2_col111[10]),
        .c_in(stage2_col111[11]),
        .s(fa_s2_c111_n360_s),
        .c_out(fa_s2_c111_n360_c)
    );

    fa fa_s2_c111_n361 (
        .a(stage2_col111[12]),
        .b(stage2_col111[13]),
        .c_in(stage2_col111[14]),
        .s(fa_s2_c111_n361_s),
        .c_out(fa_s2_c111_n361_c)
    );

    fa fa_s2_c112_n362 (
        .a(stage2_col112[0]),
        .b(stage2_col112[1]),
        .c_in(stage2_col112[2]),
        .s(fa_s2_c112_n362_s),
        .c_out(fa_s2_c112_n362_c)
    );

    fa fa_s2_c112_n363 (
        .a(stage2_col112[3]),
        .b(stage2_col112[4]),
        .c_in(stage2_col112[5]),
        .s(fa_s2_c112_n363_s),
        .c_out(fa_s2_c112_n363_c)
    );

    fa fa_s2_c112_n364 (
        .a(stage2_col112[6]),
        .b(stage2_col112[7]),
        .c_in(stage2_col112[8]),
        .s(fa_s2_c112_n364_s),
        .c_out(fa_s2_c112_n364_c)
    );

    fa fa_s2_c112_n365 (
        .a(stage2_col112[9]),
        .b(stage2_col112[10]),
        .c_in(stage2_col112[11]),
        .s(fa_s2_c112_n365_s),
        .c_out(fa_s2_c112_n365_c)
    );

    fa fa_s2_c113_n366 (
        .a(stage2_col113[0]),
        .b(stage2_col113[1]),
        .c_in(stage2_col113[2]),
        .s(fa_s2_c113_n366_s),
        .c_out(fa_s2_c113_n366_c)
    );

    fa fa_s2_c113_n367 (
        .a(stage2_col113[3]),
        .b(stage2_col113[4]),
        .c_in(stage2_col113[5]),
        .s(fa_s2_c113_n367_s),
        .c_out(fa_s2_c113_n367_c)
    );

    fa fa_s2_c113_n368 (
        .a(stage2_col113[6]),
        .b(stage2_col113[7]),
        .c_in(stage2_col113[8]),
        .s(fa_s2_c113_n368_s),
        .c_out(fa_s2_c113_n368_c)
    );

    fa fa_s2_c113_n369 (
        .a(stage2_col113[9]),
        .b(stage2_col113[10]),
        .c_in(stage2_col113[11]),
        .s(fa_s2_c113_n369_s),
        .c_out(fa_s2_c113_n369_c)
    );

    fa fa_s2_c113_n370 (
        .a(stage2_col113[12]),
        .b(stage2_col113[13]),
        .c_in(stage2_col113[14]),
        .s(fa_s2_c113_n370_s),
        .c_out(fa_s2_c113_n370_c)
    );

    fa fa_s2_c114_n371 (
        .a(stage2_col114[0]),
        .b(stage2_col114[1]),
        .c_in(stage2_col114[2]),
        .s(fa_s2_c114_n371_s),
        .c_out(fa_s2_c114_n371_c)
    );

    fa fa_s2_c114_n372 (
        .a(stage2_col114[3]),
        .b(stage2_col114[4]),
        .c_in(stage2_col114[5]),
        .s(fa_s2_c114_n372_s),
        .c_out(fa_s2_c114_n372_c)
    );

    fa fa_s2_c114_n373 (
        .a(stage2_col114[6]),
        .b(stage2_col114[7]),
        .c_in(stage2_col114[8]),
        .s(fa_s2_c114_n373_s),
        .c_out(fa_s2_c114_n373_c)
    );

    fa fa_s2_c114_n374 (
        .a(stage2_col114[9]),
        .b(stage2_col114[10]),
        .c_in(stage2_col114[11]),
        .s(fa_s2_c114_n374_s),
        .c_out(fa_s2_c114_n374_c)
    );

    fa fa_s2_c115_n375 (
        .a(stage2_col115[0]),
        .b(stage2_col115[1]),
        .c_in(stage2_col115[2]),
        .s(fa_s2_c115_n375_s),
        .c_out(fa_s2_c115_n375_c)
    );

    fa fa_s2_c115_n376 (
        .a(stage2_col115[3]),
        .b(stage2_col115[4]),
        .c_in(stage2_col115[5]),
        .s(fa_s2_c115_n376_s),
        .c_out(fa_s2_c115_n376_c)
    );

    fa fa_s2_c115_n377 (
        .a(stage2_col115[6]),
        .b(stage2_col115[7]),
        .c_in(stage2_col115[8]),
        .s(fa_s2_c115_n377_s),
        .c_out(fa_s2_c115_n377_c)
    );

    fa fa_s2_c115_n378 (
        .a(stage2_col115[9]),
        .b(stage2_col115[10]),
        .c_in(stage2_col115[11]),
        .s(fa_s2_c115_n378_s),
        .c_out(fa_s2_c115_n378_c)
    );

    fa fa_s2_c115_n379 (
        .a(stage2_col115[12]),
        .b(stage2_col115[13]),
        .c_in(stage2_col115[14]),
        .s(fa_s2_c115_n379_s),
        .c_out(fa_s2_c115_n379_c)
    );

    fa fa_s2_c116_n380 (
        .a(stage2_col116[0]),
        .b(stage2_col116[1]),
        .c_in(stage2_col116[2]),
        .s(fa_s2_c116_n380_s),
        .c_out(fa_s2_c116_n380_c)
    );

    fa fa_s2_c116_n381 (
        .a(stage2_col116[3]),
        .b(stage2_col116[4]),
        .c_in(stage2_col116[5]),
        .s(fa_s2_c116_n381_s),
        .c_out(fa_s2_c116_n381_c)
    );

    fa fa_s2_c116_n382 (
        .a(stage2_col116[6]),
        .b(stage2_col116[7]),
        .c_in(stage2_col116[8]),
        .s(fa_s2_c116_n382_s),
        .c_out(fa_s2_c116_n382_c)
    );

    fa fa_s2_c116_n383 (
        .a(stage2_col116[9]),
        .b(stage2_col116[10]),
        .c_in(stage2_col116[11]),
        .s(fa_s2_c116_n383_s),
        .c_out(fa_s2_c116_n383_c)
    );

    fa fa_s2_c117_n384 (
        .a(stage2_col117[0]),
        .b(stage2_col117[1]),
        .c_in(stage2_col117[2]),
        .s(fa_s2_c117_n384_s),
        .c_out(fa_s2_c117_n384_c)
    );

    fa fa_s2_c117_n385 (
        .a(stage2_col117[3]),
        .b(stage2_col117[4]),
        .c_in(stage2_col117[5]),
        .s(fa_s2_c117_n385_s),
        .c_out(fa_s2_c117_n385_c)
    );

    fa fa_s2_c117_n386 (
        .a(stage2_col117[6]),
        .b(stage2_col117[7]),
        .c_in(stage2_col117[8]),
        .s(fa_s2_c117_n386_s),
        .c_out(fa_s2_c117_n386_c)
    );

    fa fa_s2_c117_n387 (
        .a(stage2_col117[9]),
        .b(stage2_col117[10]),
        .c_in(stage2_col117[11]),
        .s(fa_s2_c117_n387_s),
        .c_out(fa_s2_c117_n387_c)
    );

    fa fa_s2_c117_n388 (
        .a(stage2_col117[12]),
        .b(stage2_col117[13]),
        .c_in(stage2_col117[14]),
        .s(fa_s2_c117_n388_s),
        .c_out(fa_s2_c117_n388_c)
    );

    fa fa_s2_c118_n389 (
        .a(stage2_col118[0]),
        .b(stage2_col118[1]),
        .c_in(stage2_col118[2]),
        .s(fa_s2_c118_n389_s),
        .c_out(fa_s2_c118_n389_c)
    );

    fa fa_s2_c118_n390 (
        .a(stage2_col118[3]),
        .b(stage2_col118[4]),
        .c_in(stage2_col118[5]),
        .s(fa_s2_c118_n390_s),
        .c_out(fa_s2_c118_n390_c)
    );

    fa fa_s2_c118_n391 (
        .a(stage2_col118[6]),
        .b(stage2_col118[7]),
        .c_in(stage2_col118[8]),
        .s(fa_s2_c118_n391_s),
        .c_out(fa_s2_c118_n391_c)
    );

    fa fa_s2_c118_n392 (
        .a(stage2_col118[9]),
        .b(stage2_col118[10]),
        .c_in(stage2_col118[11]),
        .s(fa_s2_c118_n392_s),
        .c_out(fa_s2_c118_n392_c)
    );

    fa fa_s2_c119_n393 (
        .a(stage2_col119[0]),
        .b(stage2_col119[1]),
        .c_in(stage2_col119[2]),
        .s(fa_s2_c119_n393_s),
        .c_out(fa_s2_c119_n393_c)
    );

    fa fa_s2_c119_n394 (
        .a(stage2_col119[3]),
        .b(stage2_col119[4]),
        .c_in(stage2_col119[5]),
        .s(fa_s2_c119_n394_s),
        .c_out(fa_s2_c119_n394_c)
    );

    fa fa_s2_c119_n395 (
        .a(stage2_col119[6]),
        .b(stage2_col119[7]),
        .c_in(stage2_col119[8]),
        .s(fa_s2_c119_n395_s),
        .c_out(fa_s2_c119_n395_c)
    );

    fa fa_s2_c119_n396 (
        .a(stage2_col119[9]),
        .b(stage2_col119[10]),
        .c_in(stage2_col119[11]),
        .s(fa_s2_c119_n396_s),
        .c_out(fa_s2_c119_n396_c)
    );

    fa fa_s2_c119_n397 (
        .a(stage2_col119[12]),
        .b(stage2_col119[13]),
        .c_in(stage2_col119[14]),
        .s(fa_s2_c119_n397_s),
        .c_out(fa_s2_c119_n397_c)
    );

    fa fa_s2_c120_n398 (
        .a(stage2_col120[0]),
        .b(stage2_col120[1]),
        .c_in(stage2_col120[2]),
        .s(fa_s2_c120_n398_s),
        .c_out(fa_s2_c120_n398_c)
    );

    fa fa_s2_c120_n399 (
        .a(stage2_col120[3]),
        .b(stage2_col120[4]),
        .c_in(stage2_col120[5]),
        .s(fa_s2_c120_n399_s),
        .c_out(fa_s2_c120_n399_c)
    );

    fa fa_s2_c120_n400 (
        .a(stage2_col120[6]),
        .b(stage2_col120[7]),
        .c_in(stage2_col120[8]),
        .s(fa_s2_c120_n400_s),
        .c_out(fa_s2_c120_n400_c)
    );

    fa fa_s2_c120_n401 (
        .a(stage2_col120[9]),
        .b(stage2_col120[10]),
        .c_in(stage2_col120[11]),
        .s(fa_s2_c120_n401_s),
        .c_out(fa_s2_c120_n401_c)
    );

    fa fa_s2_c121_n402 (
        .a(stage2_col121[0]),
        .b(stage2_col121[1]),
        .c_in(stage2_col121[2]),
        .s(fa_s2_c121_n402_s),
        .c_out(fa_s2_c121_n402_c)
    );

    fa fa_s2_c121_n403 (
        .a(stage2_col121[3]),
        .b(stage2_col121[4]),
        .c_in(stage2_col121[5]),
        .s(fa_s2_c121_n403_s),
        .c_out(fa_s2_c121_n403_c)
    );

    fa fa_s2_c121_n404 (
        .a(stage2_col121[6]),
        .b(stage2_col121[7]),
        .c_in(stage2_col121[8]),
        .s(fa_s2_c121_n404_s),
        .c_out(fa_s2_c121_n404_c)
    );

    fa fa_s2_c121_n405 (
        .a(stage2_col121[9]),
        .b(stage2_col121[10]),
        .c_in(stage2_col121[11]),
        .s(fa_s2_c121_n405_s),
        .c_out(fa_s2_c121_n405_c)
    );

    fa fa_s2_c121_n406 (
        .a(stage2_col121[12]),
        .b(stage2_col121[13]),
        .c_in(stage2_col121[14]),
        .s(fa_s2_c121_n406_s),
        .c_out(fa_s2_c121_n406_c)
    );

    fa fa_s2_c122_n407 (
        .a(stage2_col122[0]),
        .b(stage2_col122[1]),
        .c_in(stage2_col122[2]),
        .s(fa_s2_c122_n407_s),
        .c_out(fa_s2_c122_n407_c)
    );

    fa fa_s2_c122_n408 (
        .a(stage2_col122[3]),
        .b(stage2_col122[4]),
        .c_in(stage2_col122[5]),
        .s(fa_s2_c122_n408_s),
        .c_out(fa_s2_c122_n408_c)
    );

    fa fa_s2_c122_n409 (
        .a(stage2_col122[6]),
        .b(stage2_col122[7]),
        .c_in(stage2_col122[8]),
        .s(fa_s2_c122_n409_s),
        .c_out(fa_s2_c122_n409_c)
    );

    fa fa_s2_c122_n410 (
        .a(stage2_col122[9]),
        .b(stage2_col122[10]),
        .c_in(stage2_col122[11]),
        .s(fa_s2_c122_n410_s),
        .c_out(fa_s2_c122_n410_c)
    );

    fa fa_s2_c123_n411 (
        .a(stage2_col123[0]),
        .b(stage2_col123[1]),
        .c_in(stage2_col123[2]),
        .s(fa_s2_c123_n411_s),
        .c_out(fa_s2_c123_n411_c)
    );

    fa fa_s2_c123_n412 (
        .a(stage2_col123[3]),
        .b(stage2_col123[4]),
        .c_in(stage2_col123[5]),
        .s(fa_s2_c123_n412_s),
        .c_out(fa_s2_c123_n412_c)
    );

    fa fa_s2_c123_n413 (
        .a(stage2_col123[6]),
        .b(stage2_col123[7]),
        .c_in(stage2_col123[8]),
        .s(fa_s2_c123_n413_s),
        .c_out(fa_s2_c123_n413_c)
    );

    fa fa_s2_c123_n414 (
        .a(stage2_col123[9]),
        .b(stage2_col123[10]),
        .c_in(stage2_col123[11]),
        .s(fa_s2_c123_n414_s),
        .c_out(fa_s2_c123_n414_c)
    );

    fa fa_s2_c123_n415 (
        .a(stage2_col123[12]),
        .b(stage2_col123[13]),
        .c_in(stage2_col123[14]),
        .s(fa_s2_c123_n415_s),
        .c_out(fa_s2_c123_n415_c)
    );

    fa fa_s2_c124_n416 (
        .a(stage2_col124[0]),
        .b(stage2_col124[1]),
        .c_in(stage2_col124[2]),
        .s(fa_s2_c124_n416_s),
        .c_out(fa_s2_c124_n416_c)
    );

    fa fa_s2_c124_n417 (
        .a(stage2_col124[3]),
        .b(stage2_col124[4]),
        .c_in(stage2_col124[5]),
        .s(fa_s2_c124_n417_s),
        .c_out(fa_s2_c124_n417_c)
    );

    fa fa_s2_c124_n418 (
        .a(stage2_col124[6]),
        .b(stage2_col124[7]),
        .c_in(stage2_col124[8]),
        .s(fa_s2_c124_n418_s),
        .c_out(fa_s2_c124_n418_c)
    );

    fa fa_s2_c124_n419 (
        .a(stage2_col124[9]),
        .b(stage2_col124[10]),
        .c_in(stage2_col124[11]),
        .s(fa_s2_c124_n419_s),
        .c_out(fa_s2_c124_n419_c)
    );

    fa fa_s2_c125_n420 (
        .a(stage2_col125[0]),
        .b(stage2_col125[1]),
        .c_in(stage2_col125[2]),
        .s(fa_s2_c125_n420_s),
        .c_out(fa_s2_c125_n420_c)
    );

    fa fa_s2_c125_n421 (
        .a(stage2_col125[3]),
        .b(stage2_col125[4]),
        .c_in(stage2_col125[5]),
        .s(fa_s2_c125_n421_s),
        .c_out(fa_s2_c125_n421_c)
    );

    fa fa_s2_c125_n422 (
        .a(stage2_col125[6]),
        .b(stage2_col125[7]),
        .c_in(stage2_col125[8]),
        .s(fa_s2_c125_n422_s),
        .c_out(fa_s2_c125_n422_c)
    );

    fa fa_s2_c125_n423 (
        .a(stage2_col125[9]),
        .b(stage2_col125[10]),
        .c_in(stage2_col125[11]),
        .s(fa_s2_c125_n423_s),
        .c_out(fa_s2_c125_n423_c)
    );

    fa fa_s2_c125_n424 (
        .a(stage2_col125[12]),
        .b(stage2_col125[13]),
        .c_in(stage2_col125[14]),
        .s(fa_s2_c125_n424_s),
        .c_out(fa_s2_c125_n424_c)
    );

    fa fa_s2_c126_n425 (
        .a(stage2_col126[0]),
        .b(stage2_col126[1]),
        .c_in(stage2_col126[2]),
        .s(fa_s2_c126_n425_s),
        .c_out(fa_s2_c126_n425_c)
    );

    fa fa_s2_c126_n426 (
        .a(stage2_col126[3]),
        .b(stage2_col126[4]),
        .c_in(stage2_col126[5]),
        .s(fa_s2_c126_n426_s),
        .c_out(fa_s2_c126_n426_c)
    );

    fa fa_s2_c126_n427 (
        .a(stage2_col126[6]),
        .b(stage2_col126[7]),
        .c_in(stage2_col126[8]),
        .s(fa_s2_c126_n427_s),
        .c_out(fa_s2_c126_n427_c)
    );

    fa fa_s2_c126_n428 (
        .a(stage2_col126[9]),
        .b(stage2_col126[10]),
        .c_in(stage2_col126[11]),
        .s(fa_s2_c126_n428_s),
        .c_out(fa_s2_c126_n428_c)
    );

    ha ha_s2_c2_n0 (
        .a(stage2_col2[0]),
        .b(stage2_col2[1]),
        .s(ha_s2_c2_n0_s),
        .c_out(ha_s2_c2_n0_c)
    );

    // Map to Stage 3 columns
    generate
        if (PIPE) begin : gen_stage3_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage3_col0[0] <= 1'b0;
                    stage3_col1[0] <= 1'b0;
                    stage3_col2[0] <= 1'b0;
                    stage3_col3[0] <= 1'b0;
                    stage3_col3[1] <= 1'b0;
                    stage3_col4[0] <= 1'b0;
                    stage3_col5[0] <= 1'b0;
                    stage3_col5[1] <= 1'b0;
                    stage3_col5[2] <= 1'b0;
                    stage3_col6[0] <= 1'b0;
                    stage3_col6[1] <= 1'b0;
                    stage3_col7[0] <= 1'b0;
                    stage3_col7[1] <= 1'b0;
                    stage3_col8[0] <= 1'b0;
                    stage3_col8[1] <= 1'b0;
                    stage3_col9[0] <= 1'b0;
                    stage3_col9[1] <= 1'b0;
                    stage3_col10[0] <= 1'b0;
                    stage3_col10[1] <= 1'b0;
                    stage3_col11[0] <= 1'b0;
                    stage3_col11[1] <= 1'b0;
                    stage3_col12[0] <= 1'b0;
                    stage3_col12[1] <= 1'b0;
                    stage3_col13[0] <= 1'b0;
                    stage3_col13[1] <= 1'b0;
                    stage3_col13[2] <= 1'b0;
                    stage3_col13[3] <= 1'b0;
                    stage3_col14[0] <= 1'b0;
                    stage3_col14[1] <= 1'b0;
                    stage3_col14[2] <= 1'b0;
                    stage3_col15[0] <= 1'b0;
                    stage3_col15[1] <= 1'b0;
                    stage3_col15[2] <= 1'b0;
                    stage3_col16[0] <= 1'b0;
                    stage3_col16[1] <= 1'b0;
                    stage3_col16[2] <= 1'b0;
                    stage3_col17[0] <= 1'b0;
                    stage3_col17[1] <= 1'b0;
                    stage3_col17[2] <= 1'b0;
                    stage3_col18[0] <= 1'b0;
                    stage3_col18[1] <= 1'b0;
                    stage3_col18[2] <= 1'b0;
                    stage3_col19[0] <= 1'b0;
                    stage3_col19[1] <= 1'b0;
                    stage3_col19[2] <= 1'b0;
                    stage3_col19[3] <= 1'b0;
                    stage3_col19[4] <= 1'b0;
                    stage3_col20[0] <= 1'b0;
                    stage3_col20[1] <= 1'b0;
                    stage3_col20[2] <= 1'b0;
                    stage3_col20[3] <= 1'b0;
                    stage3_col21[0] <= 1'b0;
                    stage3_col21[1] <= 1'b0;
                    stage3_col21[2] <= 1'b0;
                    stage3_col21[3] <= 1'b0;
                    stage3_col22[0] <= 1'b0;
                    stage3_col22[1] <= 1'b0;
                    stage3_col22[2] <= 1'b0;
                    stage3_col22[3] <= 1'b0;
                    stage3_col23[0] <= 1'b0;
                    stage3_col23[1] <= 1'b0;
                    stage3_col23[2] <= 1'b0;
                    stage3_col23[3] <= 1'b0;
                    stage3_col24[0] <= 1'b0;
                    stage3_col24[1] <= 1'b0;
                    stage3_col24[2] <= 1'b0;
                    stage3_col24[3] <= 1'b0;
                    stage3_col25[0] <= 1'b0;
                    stage3_col25[1] <= 1'b0;
                    stage3_col25[2] <= 1'b0;
                    stage3_col25[3] <= 1'b0;
                    stage3_col26[0] <= 1'b0;
                    stage3_col26[1] <= 1'b0;
                    stage3_col26[2] <= 1'b0;
                    stage3_col26[3] <= 1'b0;
                    stage3_col27[0] <= 1'b0;
                    stage3_col27[1] <= 1'b0;
                    stage3_col27[2] <= 1'b0;
                    stage3_col27[3] <= 1'b0;
                    stage3_col27[4] <= 1'b0;
                    stage3_col27[5] <= 1'b0;
                    stage3_col28[0] <= 1'b0;
                    stage3_col28[1] <= 1'b0;
                    stage3_col28[2] <= 1'b0;
                    stage3_col28[3] <= 1'b0;
                    stage3_col28[4] <= 1'b0;
                    stage3_col29[0] <= 1'b0;
                    stage3_col29[1] <= 1'b0;
                    stage3_col29[2] <= 1'b0;
                    stage3_col29[3] <= 1'b0;
                    stage3_col29[4] <= 1'b0;
                    stage3_col30[0] <= 1'b0;
                    stage3_col30[1] <= 1'b0;
                    stage3_col30[2] <= 1'b0;
                    stage3_col30[3] <= 1'b0;
                    stage3_col30[4] <= 1'b0;
                    stage3_col31[0] <= 1'b0;
                    stage3_col31[1] <= 1'b0;
                    stage3_col31[2] <= 1'b0;
                    stage3_col31[3] <= 1'b0;
                    stage3_col31[4] <= 1'b0;
                    stage3_col32[0] <= 1'b0;
                    stage3_col32[1] <= 1'b0;
                    stage3_col32[2] <= 1'b0;
                    stage3_col32[3] <= 1'b0;
                    stage3_col32[4] <= 1'b0;
                    stage3_col32[5] <= 1'b0;
                    stage3_col32[6] <= 1'b0;
                    stage3_col33[0] <= 1'b0;
                    stage3_col33[1] <= 1'b0;
                    stage3_col33[2] <= 1'b0;
                    stage3_col33[3] <= 1'b0;
                    stage3_col33[4] <= 1'b0;
                    stage3_col33[5] <= 1'b0;
                    stage3_col34[0] <= 1'b0;
                    stage3_col34[1] <= 1'b0;
                    stage3_col34[2] <= 1'b0;
                    stage3_col34[3] <= 1'b0;
                    stage3_col34[4] <= 1'b0;
                    stage3_col34[5] <= 1'b0;
                    stage3_col35[0] <= 1'b0;
                    stage3_col35[1] <= 1'b0;
                    stage3_col35[2] <= 1'b0;
                    stage3_col35[3] <= 1'b0;
                    stage3_col35[4] <= 1'b0;
                    stage3_col35[5] <= 1'b0;
                    stage3_col36[0] <= 1'b0;
                    stage3_col36[1] <= 1'b0;
                    stage3_col36[2] <= 1'b0;
                    stage3_col36[3] <= 1'b0;
                    stage3_col36[4] <= 1'b0;
                    stage3_col36[5] <= 1'b0;
                    stage3_col37[0] <= 1'b0;
                    stage3_col37[1] <= 1'b0;
                    stage3_col37[2] <= 1'b0;
                    stage3_col37[3] <= 1'b0;
                    stage3_col37[4] <= 1'b0;
                    stage3_col37[5] <= 1'b0;
                    stage3_col38[0] <= 1'b0;
                    stage3_col38[1] <= 1'b0;
                    stage3_col38[2] <= 1'b0;
                    stage3_col38[3] <= 1'b0;
                    stage3_col38[4] <= 1'b0;
                    stage3_col38[5] <= 1'b0;
                    stage3_col39[0] <= 1'b0;
                    stage3_col39[1] <= 1'b0;
                    stage3_col39[2] <= 1'b0;
                    stage3_col39[3] <= 1'b0;
                    stage3_col39[4] <= 1'b0;
                    stage3_col39[5] <= 1'b0;
                    stage3_col40[0] <= 1'b0;
                    stage3_col40[1] <= 1'b0;
                    stage3_col40[2] <= 1'b0;
                    stage3_col40[3] <= 1'b0;
                    stage3_col40[4] <= 1'b0;
                    stage3_col40[5] <= 1'b0;
                    stage3_col40[6] <= 1'b0;
                    stage3_col40[7] <= 1'b0;
                    stage3_col41[0] <= 1'b0;
                    stage3_col41[1] <= 1'b0;
                    stage3_col41[2] <= 1'b0;
                    stage3_col41[3] <= 1'b0;
                    stage3_col41[4] <= 1'b0;
                    stage3_col41[5] <= 1'b0;
                    stage3_col41[6] <= 1'b0;
                    stage3_col42[0] <= 1'b0;
                    stage3_col42[1] <= 1'b0;
                    stage3_col42[2] <= 1'b0;
                    stage3_col42[3] <= 1'b0;
                    stage3_col42[4] <= 1'b0;
                    stage3_col42[5] <= 1'b0;
                    stage3_col42[6] <= 1'b0;
                    stage3_col43[0] <= 1'b0;
                    stage3_col43[1] <= 1'b0;
                    stage3_col43[2] <= 1'b0;
                    stage3_col43[3] <= 1'b0;
                    stage3_col43[4] <= 1'b0;
                    stage3_col43[5] <= 1'b0;
                    stage3_col43[6] <= 1'b0;
                    stage3_col44[0] <= 1'b0;
                    stage3_col44[1] <= 1'b0;
                    stage3_col44[2] <= 1'b0;
                    stage3_col44[3] <= 1'b0;
                    stage3_col44[4] <= 1'b0;
                    stage3_col44[5] <= 1'b0;
                    stage3_col44[6] <= 1'b0;
                    stage3_col45[0] <= 1'b0;
                    stage3_col45[1] <= 1'b0;
                    stage3_col45[2] <= 1'b0;
                    stage3_col45[3] <= 1'b0;
                    stage3_col45[4] <= 1'b0;
                    stage3_col45[5] <= 1'b0;
                    stage3_col45[6] <= 1'b0;
                    stage3_col46[0] <= 1'b0;
                    stage3_col46[1] <= 1'b0;
                    stage3_col46[2] <= 1'b0;
                    stage3_col46[3] <= 1'b0;
                    stage3_col46[4] <= 1'b0;
                    stage3_col46[5] <= 1'b0;
                    stage3_col46[6] <= 1'b0;
                    stage3_col46[7] <= 1'b0;
                    stage3_col46[8] <= 1'b0;
                    stage3_col47[0] <= 1'b0;
                    stage3_col47[1] <= 1'b0;
                    stage3_col47[2] <= 1'b0;
                    stage3_col47[3] <= 1'b0;
                    stage3_col47[4] <= 1'b0;
                    stage3_col47[5] <= 1'b0;
                    stage3_col47[6] <= 1'b0;
                    stage3_col47[7] <= 1'b0;
                    stage3_col48[0] <= 1'b0;
                    stage3_col48[1] <= 1'b0;
                    stage3_col48[2] <= 1'b0;
                    stage3_col48[3] <= 1'b0;
                    stage3_col48[4] <= 1'b0;
                    stage3_col48[5] <= 1'b0;
                    stage3_col48[6] <= 1'b0;
                    stage3_col48[7] <= 1'b0;
                    stage3_col49[0] <= 1'b0;
                    stage3_col49[1] <= 1'b0;
                    stage3_col49[2] <= 1'b0;
                    stage3_col49[3] <= 1'b0;
                    stage3_col49[4] <= 1'b0;
                    stage3_col49[5] <= 1'b0;
                    stage3_col49[6] <= 1'b0;
                    stage3_col49[7] <= 1'b0;
                    stage3_col50[0] <= 1'b0;
                    stage3_col50[1] <= 1'b0;
                    stage3_col50[2] <= 1'b0;
                    stage3_col50[3] <= 1'b0;
                    stage3_col50[4] <= 1'b0;
                    stage3_col50[5] <= 1'b0;
                    stage3_col50[6] <= 1'b0;
                    stage3_col50[7] <= 1'b0;
                    stage3_col51[0] <= 1'b0;
                    stage3_col51[1] <= 1'b0;
                    stage3_col51[2] <= 1'b0;
                    stage3_col51[3] <= 1'b0;
                    stage3_col51[4] <= 1'b0;
                    stage3_col51[5] <= 1'b0;
                    stage3_col51[6] <= 1'b0;
                    stage3_col51[7] <= 1'b0;
                    stage3_col52[0] <= 1'b0;
                    stage3_col52[1] <= 1'b0;
                    stage3_col52[2] <= 1'b0;
                    stage3_col52[3] <= 1'b0;
                    stage3_col52[4] <= 1'b0;
                    stage3_col52[5] <= 1'b0;
                    stage3_col52[6] <= 1'b0;
                    stage3_col52[7] <= 1'b0;
                    stage3_col53[0] <= 1'b0;
                    stage3_col53[1] <= 1'b0;
                    stage3_col53[2] <= 1'b0;
                    stage3_col53[3] <= 1'b0;
                    stage3_col53[4] <= 1'b0;
                    stage3_col53[5] <= 1'b0;
                    stage3_col53[6] <= 1'b0;
                    stage3_col53[7] <= 1'b0;
                    stage3_col54[0] <= 1'b0;
                    stage3_col54[1] <= 1'b0;
                    stage3_col54[2] <= 1'b0;
                    stage3_col54[3] <= 1'b0;
                    stage3_col54[4] <= 1'b0;
                    stage3_col54[5] <= 1'b0;
                    stage3_col54[6] <= 1'b0;
                    stage3_col54[7] <= 1'b0;
                    stage3_col54[8] <= 1'b0;
                    stage3_col54[9] <= 1'b0;
                    stage3_col55[0] <= 1'b0;
                    stage3_col55[1] <= 1'b0;
                    stage3_col55[2] <= 1'b0;
                    stage3_col55[3] <= 1'b0;
                    stage3_col55[4] <= 1'b0;
                    stage3_col55[5] <= 1'b0;
                    stage3_col55[6] <= 1'b0;
                    stage3_col55[7] <= 1'b0;
                    stage3_col55[8] <= 1'b0;
                    stage3_col56[0] <= 1'b0;
                    stage3_col56[1] <= 1'b0;
                    stage3_col56[2] <= 1'b0;
                    stage3_col56[3] <= 1'b0;
                    stage3_col56[4] <= 1'b0;
                    stage3_col56[5] <= 1'b0;
                    stage3_col56[6] <= 1'b0;
                    stage3_col56[7] <= 1'b0;
                    stage3_col56[8] <= 1'b0;
                    stage3_col57[0] <= 1'b0;
                    stage3_col57[1] <= 1'b0;
                    stage3_col57[2] <= 1'b0;
                    stage3_col57[3] <= 1'b0;
                    stage3_col57[4] <= 1'b0;
                    stage3_col57[5] <= 1'b0;
                    stage3_col57[6] <= 1'b0;
                    stage3_col57[7] <= 1'b0;
                    stage3_col57[8] <= 1'b0;
                    stage3_col58[0] <= 1'b0;
                    stage3_col58[1] <= 1'b0;
                    stage3_col58[2] <= 1'b0;
                    stage3_col58[3] <= 1'b0;
                    stage3_col58[4] <= 1'b0;
                    stage3_col58[5] <= 1'b0;
                    stage3_col58[6] <= 1'b0;
                    stage3_col58[7] <= 1'b0;
                    stage3_col58[8] <= 1'b0;
                    stage3_col59[0] <= 1'b0;
                    stage3_col59[1] <= 1'b0;
                    stage3_col59[2] <= 1'b0;
                    stage3_col59[3] <= 1'b0;
                    stage3_col59[4] <= 1'b0;
                    stage3_col59[5] <= 1'b0;
                    stage3_col59[6] <= 1'b0;
                    stage3_col59[7] <= 1'b0;
                    stage3_col59[8] <= 1'b0;
                    stage3_col59[9] <= 1'b0;
                    stage3_col59[10] <= 1'b0;
                    stage3_col60[0] <= 1'b0;
                    stage3_col60[1] <= 1'b0;
                    stage3_col60[2] <= 1'b0;
                    stage3_col60[3] <= 1'b0;
                    stage3_col60[4] <= 1'b0;
                    stage3_col60[5] <= 1'b0;
                    stage3_col60[6] <= 1'b0;
                    stage3_col60[7] <= 1'b0;
                    stage3_col60[8] <= 1'b0;
                    stage3_col60[9] <= 1'b0;
                    stage3_col61[0] <= 1'b0;
                    stage3_col61[1] <= 1'b0;
                    stage3_col61[2] <= 1'b0;
                    stage3_col61[3] <= 1'b0;
                    stage3_col61[4] <= 1'b0;
                    stage3_col61[5] <= 1'b0;
                    stage3_col61[6] <= 1'b0;
                    stage3_col61[7] <= 1'b0;
                    stage3_col61[8] <= 1'b0;
                    stage3_col61[9] <= 1'b0;
                    stage3_col62[0] <= 1'b0;
                    stage3_col62[1] <= 1'b0;
                    stage3_col62[2] <= 1'b0;
                    stage3_col62[3] <= 1'b0;
                    stage3_col62[4] <= 1'b0;
                    stage3_col62[5] <= 1'b0;
                    stage3_col62[6] <= 1'b0;
                    stage3_col62[7] <= 1'b0;
                    stage3_col62[8] <= 1'b0;
                    stage3_col62[9] <= 1'b0;
                    stage3_col63[0] <= 1'b0;
                    stage3_col63[1] <= 1'b0;
                    stage3_col63[2] <= 1'b0;
                    stage3_col63[3] <= 1'b0;
                    stage3_col63[4] <= 1'b0;
                    stage3_col63[5] <= 1'b0;
                    stage3_col63[6] <= 1'b0;
                    stage3_col63[7] <= 1'b0;
                    stage3_col63[8] <= 1'b0;
                    stage3_col63[9] <= 1'b0;
                    stage3_col64[0] <= 1'b0;
                    stage3_col64[1] <= 1'b0;
                    stage3_col64[2] <= 1'b0;
                    stage3_col64[3] <= 1'b0;
                    stage3_col64[4] <= 1'b0;
                    stage3_col64[5] <= 1'b0;
                    stage3_col64[6] <= 1'b0;
                    stage3_col64[7] <= 1'b0;
                    stage3_col64[8] <= 1'b0;
                    stage3_col64[9] <= 1'b0;
                    stage3_col64[10] <= 1'b0;
                    stage3_col65[0] <= 1'b0;
                    stage3_col65[1] <= 1'b0;
                    stage3_col65[2] <= 1'b0;
                    stage3_col65[3] <= 1'b0;
                    stage3_col65[4] <= 1'b0;
                    stage3_col65[5] <= 1'b0;
                    stage3_col65[6] <= 1'b0;
                    stage3_col65[7] <= 1'b0;
                    stage3_col65[8] <= 1'b0;
                    stage3_col65[9] <= 1'b0;
                    stage3_col66[0] <= 1'b0;
                    stage3_col66[1] <= 1'b0;
                    stage3_col66[2] <= 1'b0;
                    stage3_col66[3] <= 1'b0;
                    stage3_col66[4] <= 1'b0;
                    stage3_col66[5] <= 1'b0;
                    stage3_col66[6] <= 1'b0;
                    stage3_col66[7] <= 1'b0;
                    stage3_col66[8] <= 1'b0;
                    stage3_col66[9] <= 1'b0;
                    stage3_col66[10] <= 1'b0;
                    stage3_col67[0] <= 1'b0;
                    stage3_col67[1] <= 1'b0;
                    stage3_col67[2] <= 1'b0;
                    stage3_col67[3] <= 1'b0;
                    stage3_col67[4] <= 1'b0;
                    stage3_col67[5] <= 1'b0;
                    stage3_col67[6] <= 1'b0;
                    stage3_col67[7] <= 1'b0;
                    stage3_col67[8] <= 1'b0;
                    stage3_col67[9] <= 1'b0;
                    stage3_col68[0] <= 1'b0;
                    stage3_col68[1] <= 1'b0;
                    stage3_col68[2] <= 1'b0;
                    stage3_col68[3] <= 1'b0;
                    stage3_col68[4] <= 1'b0;
                    stage3_col68[5] <= 1'b0;
                    stage3_col68[6] <= 1'b0;
                    stage3_col68[7] <= 1'b0;
                    stage3_col68[8] <= 1'b0;
                    stage3_col68[9] <= 1'b0;
                    stage3_col68[10] <= 1'b0;
                    stage3_col69[0] <= 1'b0;
                    stage3_col69[1] <= 1'b0;
                    stage3_col69[2] <= 1'b0;
                    stage3_col69[3] <= 1'b0;
                    stage3_col69[4] <= 1'b0;
                    stage3_col69[5] <= 1'b0;
                    stage3_col69[6] <= 1'b0;
                    stage3_col69[7] <= 1'b0;
                    stage3_col69[8] <= 1'b0;
                    stage3_col69[9] <= 1'b0;
                    stage3_col70[0] <= 1'b0;
                    stage3_col70[1] <= 1'b0;
                    stage3_col70[2] <= 1'b0;
                    stage3_col70[3] <= 1'b0;
                    stage3_col70[4] <= 1'b0;
                    stage3_col70[5] <= 1'b0;
                    stage3_col70[6] <= 1'b0;
                    stage3_col70[7] <= 1'b0;
                    stage3_col70[8] <= 1'b0;
                    stage3_col70[9] <= 1'b0;
                    stage3_col70[10] <= 1'b0;
                    stage3_col71[0] <= 1'b0;
                    stage3_col71[1] <= 1'b0;
                    stage3_col71[2] <= 1'b0;
                    stage3_col71[3] <= 1'b0;
                    stage3_col71[4] <= 1'b0;
                    stage3_col71[5] <= 1'b0;
                    stage3_col71[6] <= 1'b0;
                    stage3_col71[7] <= 1'b0;
                    stage3_col71[8] <= 1'b0;
                    stage3_col71[9] <= 1'b0;
                    stage3_col72[0] <= 1'b0;
                    stage3_col72[1] <= 1'b0;
                    stage3_col72[2] <= 1'b0;
                    stage3_col72[3] <= 1'b0;
                    stage3_col72[4] <= 1'b0;
                    stage3_col72[5] <= 1'b0;
                    stage3_col72[6] <= 1'b0;
                    stage3_col72[7] <= 1'b0;
                    stage3_col72[8] <= 1'b0;
                    stage3_col72[9] <= 1'b0;
                    stage3_col72[10] <= 1'b0;
                    stage3_col73[0] <= 1'b0;
                    stage3_col73[1] <= 1'b0;
                    stage3_col73[2] <= 1'b0;
                    stage3_col73[3] <= 1'b0;
                    stage3_col73[4] <= 1'b0;
                    stage3_col73[5] <= 1'b0;
                    stage3_col73[6] <= 1'b0;
                    stage3_col73[7] <= 1'b0;
                    stage3_col73[8] <= 1'b0;
                    stage3_col73[9] <= 1'b0;
                    stage3_col74[0] <= 1'b0;
                    stage3_col74[1] <= 1'b0;
                    stage3_col74[2] <= 1'b0;
                    stage3_col74[3] <= 1'b0;
                    stage3_col74[4] <= 1'b0;
                    stage3_col74[5] <= 1'b0;
                    stage3_col74[6] <= 1'b0;
                    stage3_col74[7] <= 1'b0;
                    stage3_col74[8] <= 1'b0;
                    stage3_col74[9] <= 1'b0;
                    stage3_col74[10] <= 1'b0;
                    stage3_col75[0] <= 1'b0;
                    stage3_col75[1] <= 1'b0;
                    stage3_col75[2] <= 1'b0;
                    stage3_col75[3] <= 1'b0;
                    stage3_col75[4] <= 1'b0;
                    stage3_col75[5] <= 1'b0;
                    stage3_col75[6] <= 1'b0;
                    stage3_col75[7] <= 1'b0;
                    stage3_col75[8] <= 1'b0;
                    stage3_col75[9] <= 1'b0;
                    stage3_col76[0] <= 1'b0;
                    stage3_col76[1] <= 1'b0;
                    stage3_col76[2] <= 1'b0;
                    stage3_col76[3] <= 1'b0;
                    stage3_col76[4] <= 1'b0;
                    stage3_col76[5] <= 1'b0;
                    stage3_col76[6] <= 1'b0;
                    stage3_col76[7] <= 1'b0;
                    stage3_col76[8] <= 1'b0;
                    stage3_col76[9] <= 1'b0;
                    stage3_col76[10] <= 1'b0;
                    stage3_col77[0] <= 1'b0;
                    stage3_col77[1] <= 1'b0;
                    stage3_col77[2] <= 1'b0;
                    stage3_col77[3] <= 1'b0;
                    stage3_col77[4] <= 1'b0;
                    stage3_col77[5] <= 1'b0;
                    stage3_col77[6] <= 1'b0;
                    stage3_col77[7] <= 1'b0;
                    stage3_col77[8] <= 1'b0;
                    stage3_col77[9] <= 1'b0;
                    stage3_col78[0] <= 1'b0;
                    stage3_col78[1] <= 1'b0;
                    stage3_col78[2] <= 1'b0;
                    stage3_col78[3] <= 1'b0;
                    stage3_col78[4] <= 1'b0;
                    stage3_col78[5] <= 1'b0;
                    stage3_col78[6] <= 1'b0;
                    stage3_col78[7] <= 1'b0;
                    stage3_col78[8] <= 1'b0;
                    stage3_col78[9] <= 1'b0;
                    stage3_col78[10] <= 1'b0;
                    stage3_col79[0] <= 1'b0;
                    stage3_col79[1] <= 1'b0;
                    stage3_col79[2] <= 1'b0;
                    stage3_col79[3] <= 1'b0;
                    stage3_col79[4] <= 1'b0;
                    stage3_col79[5] <= 1'b0;
                    stage3_col79[6] <= 1'b0;
                    stage3_col79[7] <= 1'b0;
                    stage3_col79[8] <= 1'b0;
                    stage3_col79[9] <= 1'b0;
                    stage3_col80[0] <= 1'b0;
                    stage3_col80[1] <= 1'b0;
                    stage3_col80[2] <= 1'b0;
                    stage3_col80[3] <= 1'b0;
                    stage3_col80[4] <= 1'b0;
                    stage3_col80[5] <= 1'b0;
                    stage3_col80[6] <= 1'b0;
                    stage3_col80[7] <= 1'b0;
                    stage3_col80[8] <= 1'b0;
                    stage3_col80[9] <= 1'b0;
                    stage3_col80[10] <= 1'b0;
                    stage3_col81[0] <= 1'b0;
                    stage3_col81[1] <= 1'b0;
                    stage3_col81[2] <= 1'b0;
                    stage3_col81[3] <= 1'b0;
                    stage3_col81[4] <= 1'b0;
                    stage3_col81[5] <= 1'b0;
                    stage3_col81[6] <= 1'b0;
                    stage3_col81[7] <= 1'b0;
                    stage3_col81[8] <= 1'b0;
                    stage3_col81[9] <= 1'b0;
                    stage3_col82[0] <= 1'b0;
                    stage3_col82[1] <= 1'b0;
                    stage3_col82[2] <= 1'b0;
                    stage3_col82[3] <= 1'b0;
                    stage3_col82[4] <= 1'b0;
                    stage3_col82[5] <= 1'b0;
                    stage3_col82[6] <= 1'b0;
                    stage3_col82[7] <= 1'b0;
                    stage3_col82[8] <= 1'b0;
                    stage3_col82[9] <= 1'b0;
                    stage3_col82[10] <= 1'b0;
                    stage3_col83[0] <= 1'b0;
                    stage3_col83[1] <= 1'b0;
                    stage3_col83[2] <= 1'b0;
                    stage3_col83[3] <= 1'b0;
                    stage3_col83[4] <= 1'b0;
                    stage3_col83[5] <= 1'b0;
                    stage3_col83[6] <= 1'b0;
                    stage3_col83[7] <= 1'b0;
                    stage3_col83[8] <= 1'b0;
                    stage3_col83[9] <= 1'b0;
                    stage3_col84[0] <= 1'b0;
                    stage3_col84[1] <= 1'b0;
                    stage3_col84[2] <= 1'b0;
                    stage3_col84[3] <= 1'b0;
                    stage3_col84[4] <= 1'b0;
                    stage3_col84[5] <= 1'b0;
                    stage3_col84[6] <= 1'b0;
                    stage3_col84[7] <= 1'b0;
                    stage3_col84[8] <= 1'b0;
                    stage3_col84[9] <= 1'b0;
                    stage3_col84[10] <= 1'b0;
                    stage3_col85[0] <= 1'b0;
                    stage3_col85[1] <= 1'b0;
                    stage3_col85[2] <= 1'b0;
                    stage3_col85[3] <= 1'b0;
                    stage3_col85[4] <= 1'b0;
                    stage3_col85[5] <= 1'b0;
                    stage3_col85[6] <= 1'b0;
                    stage3_col85[7] <= 1'b0;
                    stage3_col85[8] <= 1'b0;
                    stage3_col85[9] <= 1'b0;
                    stage3_col86[0] <= 1'b0;
                    stage3_col86[1] <= 1'b0;
                    stage3_col86[2] <= 1'b0;
                    stage3_col86[3] <= 1'b0;
                    stage3_col86[4] <= 1'b0;
                    stage3_col86[5] <= 1'b0;
                    stage3_col86[6] <= 1'b0;
                    stage3_col86[7] <= 1'b0;
                    stage3_col86[8] <= 1'b0;
                    stage3_col86[9] <= 1'b0;
                    stage3_col86[10] <= 1'b0;
                    stage3_col87[0] <= 1'b0;
                    stage3_col87[1] <= 1'b0;
                    stage3_col87[2] <= 1'b0;
                    stage3_col87[3] <= 1'b0;
                    stage3_col87[4] <= 1'b0;
                    stage3_col87[5] <= 1'b0;
                    stage3_col87[6] <= 1'b0;
                    stage3_col87[7] <= 1'b0;
                    stage3_col87[8] <= 1'b0;
                    stage3_col87[9] <= 1'b0;
                    stage3_col88[0] <= 1'b0;
                    stage3_col88[1] <= 1'b0;
                    stage3_col88[2] <= 1'b0;
                    stage3_col88[3] <= 1'b0;
                    stage3_col88[4] <= 1'b0;
                    stage3_col88[5] <= 1'b0;
                    stage3_col88[6] <= 1'b0;
                    stage3_col88[7] <= 1'b0;
                    stage3_col88[8] <= 1'b0;
                    stage3_col88[9] <= 1'b0;
                    stage3_col88[10] <= 1'b0;
                    stage3_col89[0] <= 1'b0;
                    stage3_col89[1] <= 1'b0;
                    stage3_col89[2] <= 1'b0;
                    stage3_col89[3] <= 1'b0;
                    stage3_col89[4] <= 1'b0;
                    stage3_col89[5] <= 1'b0;
                    stage3_col89[6] <= 1'b0;
                    stage3_col89[7] <= 1'b0;
                    stage3_col89[8] <= 1'b0;
                    stage3_col89[9] <= 1'b0;
                    stage3_col90[0] <= 1'b0;
                    stage3_col90[1] <= 1'b0;
                    stage3_col90[2] <= 1'b0;
                    stage3_col90[3] <= 1'b0;
                    stage3_col90[4] <= 1'b0;
                    stage3_col90[5] <= 1'b0;
                    stage3_col90[6] <= 1'b0;
                    stage3_col90[7] <= 1'b0;
                    stage3_col90[8] <= 1'b0;
                    stage3_col90[9] <= 1'b0;
                    stage3_col90[10] <= 1'b0;
                    stage3_col91[0] <= 1'b0;
                    stage3_col91[1] <= 1'b0;
                    stage3_col91[2] <= 1'b0;
                    stage3_col91[3] <= 1'b0;
                    stage3_col91[4] <= 1'b0;
                    stage3_col91[5] <= 1'b0;
                    stage3_col91[6] <= 1'b0;
                    stage3_col91[7] <= 1'b0;
                    stage3_col91[8] <= 1'b0;
                    stage3_col91[9] <= 1'b0;
                    stage3_col92[0] <= 1'b0;
                    stage3_col92[1] <= 1'b0;
                    stage3_col92[2] <= 1'b0;
                    stage3_col92[3] <= 1'b0;
                    stage3_col92[4] <= 1'b0;
                    stage3_col92[5] <= 1'b0;
                    stage3_col92[6] <= 1'b0;
                    stage3_col92[7] <= 1'b0;
                    stage3_col92[8] <= 1'b0;
                    stage3_col92[9] <= 1'b0;
                    stage3_col92[10] <= 1'b0;
                    stage3_col93[0] <= 1'b0;
                    stage3_col93[1] <= 1'b0;
                    stage3_col93[2] <= 1'b0;
                    stage3_col93[3] <= 1'b0;
                    stage3_col93[4] <= 1'b0;
                    stage3_col93[5] <= 1'b0;
                    stage3_col93[6] <= 1'b0;
                    stage3_col93[7] <= 1'b0;
                    stage3_col93[8] <= 1'b0;
                    stage3_col93[9] <= 1'b0;
                    stage3_col94[0] <= 1'b0;
                    stage3_col94[1] <= 1'b0;
                    stage3_col94[2] <= 1'b0;
                    stage3_col94[3] <= 1'b0;
                    stage3_col94[4] <= 1'b0;
                    stage3_col94[5] <= 1'b0;
                    stage3_col94[6] <= 1'b0;
                    stage3_col94[7] <= 1'b0;
                    stage3_col94[8] <= 1'b0;
                    stage3_col94[9] <= 1'b0;
                    stage3_col94[10] <= 1'b0;
                    stage3_col95[0] <= 1'b0;
                    stage3_col95[1] <= 1'b0;
                    stage3_col95[2] <= 1'b0;
                    stage3_col95[3] <= 1'b0;
                    stage3_col95[4] <= 1'b0;
                    stage3_col95[5] <= 1'b0;
                    stage3_col95[6] <= 1'b0;
                    stage3_col95[7] <= 1'b0;
                    stage3_col95[8] <= 1'b0;
                    stage3_col95[9] <= 1'b0;
                    stage3_col96[0] <= 1'b0;
                    stage3_col96[1] <= 1'b0;
                    stage3_col96[2] <= 1'b0;
                    stage3_col96[3] <= 1'b0;
                    stage3_col96[4] <= 1'b0;
                    stage3_col96[5] <= 1'b0;
                    stage3_col96[6] <= 1'b0;
                    stage3_col96[7] <= 1'b0;
                    stage3_col96[8] <= 1'b0;
                    stage3_col96[9] <= 1'b0;
                    stage3_col96[10] <= 1'b0;
                    stage3_col97[0] <= 1'b0;
                    stage3_col97[1] <= 1'b0;
                    stage3_col97[2] <= 1'b0;
                    stage3_col97[3] <= 1'b0;
                    stage3_col97[4] <= 1'b0;
                    stage3_col97[5] <= 1'b0;
                    stage3_col97[6] <= 1'b0;
                    stage3_col97[7] <= 1'b0;
                    stage3_col97[8] <= 1'b0;
                    stage3_col97[9] <= 1'b0;
                    stage3_col98[0] <= 1'b0;
                    stage3_col98[1] <= 1'b0;
                    stage3_col98[2] <= 1'b0;
                    stage3_col98[3] <= 1'b0;
                    stage3_col98[4] <= 1'b0;
                    stage3_col98[5] <= 1'b0;
                    stage3_col98[6] <= 1'b0;
                    stage3_col98[7] <= 1'b0;
                    stage3_col98[8] <= 1'b0;
                    stage3_col98[9] <= 1'b0;
                    stage3_col98[10] <= 1'b0;
                    stage3_col99[0] <= 1'b0;
                    stage3_col99[1] <= 1'b0;
                    stage3_col99[2] <= 1'b0;
                    stage3_col99[3] <= 1'b0;
                    stage3_col99[4] <= 1'b0;
                    stage3_col99[5] <= 1'b0;
                    stage3_col99[6] <= 1'b0;
                    stage3_col99[7] <= 1'b0;
                    stage3_col99[8] <= 1'b0;
                    stage3_col99[9] <= 1'b0;
                    stage3_col100[0] <= 1'b0;
                    stage3_col100[1] <= 1'b0;
                    stage3_col100[2] <= 1'b0;
                    stage3_col100[3] <= 1'b0;
                    stage3_col100[4] <= 1'b0;
                    stage3_col100[5] <= 1'b0;
                    stage3_col100[6] <= 1'b0;
                    stage3_col100[7] <= 1'b0;
                    stage3_col100[8] <= 1'b0;
                    stage3_col100[9] <= 1'b0;
                    stage3_col100[10] <= 1'b0;
                    stage3_col101[0] <= 1'b0;
                    stage3_col101[1] <= 1'b0;
                    stage3_col101[2] <= 1'b0;
                    stage3_col101[3] <= 1'b0;
                    stage3_col101[4] <= 1'b0;
                    stage3_col101[5] <= 1'b0;
                    stage3_col101[6] <= 1'b0;
                    stage3_col101[7] <= 1'b0;
                    stage3_col101[8] <= 1'b0;
                    stage3_col101[9] <= 1'b0;
                    stage3_col102[0] <= 1'b0;
                    stage3_col102[1] <= 1'b0;
                    stage3_col102[2] <= 1'b0;
                    stage3_col102[3] <= 1'b0;
                    stage3_col102[4] <= 1'b0;
                    stage3_col102[5] <= 1'b0;
                    stage3_col102[6] <= 1'b0;
                    stage3_col102[7] <= 1'b0;
                    stage3_col102[8] <= 1'b0;
                    stage3_col102[9] <= 1'b0;
                    stage3_col102[10] <= 1'b0;
                    stage3_col103[0] <= 1'b0;
                    stage3_col103[1] <= 1'b0;
                    stage3_col103[2] <= 1'b0;
                    stage3_col103[3] <= 1'b0;
                    stage3_col103[4] <= 1'b0;
                    stage3_col103[5] <= 1'b0;
                    stage3_col103[6] <= 1'b0;
                    stage3_col103[7] <= 1'b0;
                    stage3_col103[8] <= 1'b0;
                    stage3_col103[9] <= 1'b0;
                    stage3_col104[0] <= 1'b0;
                    stage3_col104[1] <= 1'b0;
                    stage3_col104[2] <= 1'b0;
                    stage3_col104[3] <= 1'b0;
                    stage3_col104[4] <= 1'b0;
                    stage3_col104[5] <= 1'b0;
                    stage3_col104[6] <= 1'b0;
                    stage3_col104[7] <= 1'b0;
                    stage3_col104[8] <= 1'b0;
                    stage3_col104[9] <= 1'b0;
                    stage3_col104[10] <= 1'b0;
                    stage3_col105[0] <= 1'b0;
                    stage3_col105[1] <= 1'b0;
                    stage3_col105[2] <= 1'b0;
                    stage3_col105[3] <= 1'b0;
                    stage3_col105[4] <= 1'b0;
                    stage3_col105[5] <= 1'b0;
                    stage3_col105[6] <= 1'b0;
                    stage3_col105[7] <= 1'b0;
                    stage3_col105[8] <= 1'b0;
                    stage3_col105[9] <= 1'b0;
                    stage3_col106[0] <= 1'b0;
                    stage3_col106[1] <= 1'b0;
                    stage3_col106[2] <= 1'b0;
                    stage3_col106[3] <= 1'b0;
                    stage3_col106[4] <= 1'b0;
                    stage3_col106[5] <= 1'b0;
                    stage3_col106[6] <= 1'b0;
                    stage3_col106[7] <= 1'b0;
                    stage3_col106[8] <= 1'b0;
                    stage3_col106[9] <= 1'b0;
                    stage3_col106[10] <= 1'b0;
                    stage3_col107[0] <= 1'b0;
                    stage3_col107[1] <= 1'b0;
                    stage3_col107[2] <= 1'b0;
                    stage3_col107[3] <= 1'b0;
                    stage3_col107[4] <= 1'b0;
                    stage3_col107[5] <= 1'b0;
                    stage3_col107[6] <= 1'b0;
                    stage3_col107[7] <= 1'b0;
                    stage3_col107[8] <= 1'b0;
                    stage3_col107[9] <= 1'b0;
                    stage3_col108[0] <= 1'b0;
                    stage3_col108[1] <= 1'b0;
                    stage3_col108[2] <= 1'b0;
                    stage3_col108[3] <= 1'b0;
                    stage3_col108[4] <= 1'b0;
                    stage3_col108[5] <= 1'b0;
                    stage3_col108[6] <= 1'b0;
                    stage3_col108[7] <= 1'b0;
                    stage3_col108[8] <= 1'b0;
                    stage3_col108[9] <= 1'b0;
                    stage3_col108[10] <= 1'b0;
                    stage3_col109[0] <= 1'b0;
                    stage3_col109[1] <= 1'b0;
                    stage3_col109[2] <= 1'b0;
                    stage3_col109[3] <= 1'b0;
                    stage3_col109[4] <= 1'b0;
                    stage3_col109[5] <= 1'b0;
                    stage3_col109[6] <= 1'b0;
                    stage3_col109[7] <= 1'b0;
                    stage3_col109[8] <= 1'b0;
                    stage3_col109[9] <= 1'b0;
                    stage3_col110[0] <= 1'b0;
                    stage3_col110[1] <= 1'b0;
                    stage3_col110[2] <= 1'b0;
                    stage3_col110[3] <= 1'b0;
                    stage3_col110[4] <= 1'b0;
                    stage3_col110[5] <= 1'b0;
                    stage3_col110[6] <= 1'b0;
                    stage3_col110[7] <= 1'b0;
                    stage3_col110[8] <= 1'b0;
                    stage3_col110[9] <= 1'b0;
                    stage3_col110[10] <= 1'b0;
                    stage3_col111[0] <= 1'b0;
                    stage3_col111[1] <= 1'b0;
                    stage3_col111[2] <= 1'b0;
                    stage3_col111[3] <= 1'b0;
                    stage3_col111[4] <= 1'b0;
                    stage3_col111[5] <= 1'b0;
                    stage3_col111[6] <= 1'b0;
                    stage3_col111[7] <= 1'b0;
                    stage3_col111[8] <= 1'b0;
                    stage3_col111[9] <= 1'b0;
                    stage3_col112[0] <= 1'b0;
                    stage3_col112[1] <= 1'b0;
                    stage3_col112[2] <= 1'b0;
                    stage3_col112[3] <= 1'b0;
                    stage3_col112[4] <= 1'b0;
                    stage3_col112[5] <= 1'b0;
                    stage3_col112[6] <= 1'b0;
                    stage3_col112[7] <= 1'b0;
                    stage3_col112[8] <= 1'b0;
                    stage3_col112[9] <= 1'b0;
                    stage3_col112[10] <= 1'b0;
                    stage3_col113[0] <= 1'b0;
                    stage3_col113[1] <= 1'b0;
                    stage3_col113[2] <= 1'b0;
                    stage3_col113[3] <= 1'b0;
                    stage3_col113[4] <= 1'b0;
                    stage3_col113[5] <= 1'b0;
                    stage3_col113[6] <= 1'b0;
                    stage3_col113[7] <= 1'b0;
                    stage3_col113[8] <= 1'b0;
                    stage3_col113[9] <= 1'b0;
                    stage3_col114[0] <= 1'b0;
                    stage3_col114[1] <= 1'b0;
                    stage3_col114[2] <= 1'b0;
                    stage3_col114[3] <= 1'b0;
                    stage3_col114[4] <= 1'b0;
                    stage3_col114[5] <= 1'b0;
                    stage3_col114[6] <= 1'b0;
                    stage3_col114[7] <= 1'b0;
                    stage3_col114[8] <= 1'b0;
                    stage3_col114[9] <= 1'b0;
                    stage3_col114[10] <= 1'b0;
                    stage3_col115[0] <= 1'b0;
                    stage3_col115[1] <= 1'b0;
                    stage3_col115[2] <= 1'b0;
                    stage3_col115[3] <= 1'b0;
                    stage3_col115[4] <= 1'b0;
                    stage3_col115[5] <= 1'b0;
                    stage3_col115[6] <= 1'b0;
                    stage3_col115[7] <= 1'b0;
                    stage3_col115[8] <= 1'b0;
                    stage3_col115[9] <= 1'b0;
                    stage3_col116[0] <= 1'b0;
                    stage3_col116[1] <= 1'b0;
                    stage3_col116[2] <= 1'b0;
                    stage3_col116[3] <= 1'b0;
                    stage3_col116[4] <= 1'b0;
                    stage3_col116[5] <= 1'b0;
                    stage3_col116[6] <= 1'b0;
                    stage3_col116[7] <= 1'b0;
                    stage3_col116[8] <= 1'b0;
                    stage3_col116[9] <= 1'b0;
                    stage3_col116[10] <= 1'b0;
                    stage3_col117[0] <= 1'b0;
                    stage3_col117[1] <= 1'b0;
                    stage3_col117[2] <= 1'b0;
                    stage3_col117[3] <= 1'b0;
                    stage3_col117[4] <= 1'b0;
                    stage3_col117[5] <= 1'b0;
                    stage3_col117[6] <= 1'b0;
                    stage3_col117[7] <= 1'b0;
                    stage3_col117[8] <= 1'b0;
                    stage3_col117[9] <= 1'b0;
                    stage3_col118[0] <= 1'b0;
                    stage3_col118[1] <= 1'b0;
                    stage3_col118[2] <= 1'b0;
                    stage3_col118[3] <= 1'b0;
                    stage3_col118[4] <= 1'b0;
                    stage3_col118[5] <= 1'b0;
                    stage3_col118[6] <= 1'b0;
                    stage3_col118[7] <= 1'b0;
                    stage3_col118[8] <= 1'b0;
                    stage3_col118[9] <= 1'b0;
                    stage3_col118[10] <= 1'b0;
                    stage3_col119[0] <= 1'b0;
                    stage3_col119[1] <= 1'b0;
                    stage3_col119[2] <= 1'b0;
                    stage3_col119[3] <= 1'b0;
                    stage3_col119[4] <= 1'b0;
                    stage3_col119[5] <= 1'b0;
                    stage3_col119[6] <= 1'b0;
                    stage3_col119[7] <= 1'b0;
                    stage3_col119[8] <= 1'b0;
                    stage3_col119[9] <= 1'b0;
                    stage3_col120[0] <= 1'b0;
                    stage3_col120[1] <= 1'b0;
                    stage3_col120[2] <= 1'b0;
                    stage3_col120[3] <= 1'b0;
                    stage3_col120[4] <= 1'b0;
                    stage3_col120[5] <= 1'b0;
                    stage3_col120[6] <= 1'b0;
                    stage3_col120[7] <= 1'b0;
                    stage3_col120[8] <= 1'b0;
                    stage3_col120[9] <= 1'b0;
                    stage3_col120[10] <= 1'b0;
                    stage3_col121[0] <= 1'b0;
                    stage3_col121[1] <= 1'b0;
                    stage3_col121[2] <= 1'b0;
                    stage3_col121[3] <= 1'b0;
                    stage3_col121[4] <= 1'b0;
                    stage3_col121[5] <= 1'b0;
                    stage3_col121[6] <= 1'b0;
                    stage3_col121[7] <= 1'b0;
                    stage3_col121[8] <= 1'b0;
                    stage3_col121[9] <= 1'b0;
                    stage3_col122[0] <= 1'b0;
                    stage3_col122[1] <= 1'b0;
                    stage3_col122[2] <= 1'b0;
                    stage3_col122[3] <= 1'b0;
                    stage3_col122[4] <= 1'b0;
                    stage3_col122[5] <= 1'b0;
                    stage3_col122[6] <= 1'b0;
                    stage3_col122[7] <= 1'b0;
                    stage3_col122[8] <= 1'b0;
                    stage3_col122[9] <= 1'b0;
                    stage3_col122[10] <= 1'b0;
                    stage3_col123[0] <= 1'b0;
                    stage3_col123[1] <= 1'b0;
                    stage3_col123[2] <= 1'b0;
                    stage3_col123[3] <= 1'b0;
                    stage3_col123[4] <= 1'b0;
                    stage3_col123[5] <= 1'b0;
                    stage3_col123[6] <= 1'b0;
                    stage3_col123[7] <= 1'b0;
                    stage3_col123[8] <= 1'b0;
                    stage3_col123[9] <= 1'b0;
                    stage3_col124[0] <= 1'b0;
                    stage3_col124[1] <= 1'b0;
                    stage3_col124[2] <= 1'b0;
                    stage3_col124[3] <= 1'b0;
                    stage3_col124[4] <= 1'b0;
                    stage3_col124[5] <= 1'b0;
                    stage3_col124[6] <= 1'b0;
                    stage3_col124[7] <= 1'b0;
                    stage3_col124[8] <= 1'b0;
                    stage3_col124[9] <= 1'b0;
                    stage3_col124[10] <= 1'b0;
                    stage3_col125[0] <= 1'b0;
                    stage3_col125[1] <= 1'b0;
                    stage3_col125[2] <= 1'b0;
                    stage3_col125[3] <= 1'b0;
                    stage3_col125[4] <= 1'b0;
                    stage3_col125[5] <= 1'b0;
                    stage3_col125[6] <= 1'b0;
                    stage3_col125[7] <= 1'b0;
                    stage3_col125[8] <= 1'b0;
                    stage3_col125[9] <= 1'b0;
                    stage3_col126[0] <= 1'b0;
                    stage3_col126[1] <= 1'b0;
                    stage3_col126[2] <= 1'b0;
                    stage3_col126[3] <= 1'b0;
                    stage3_col126[4] <= 1'b0;
                    stage3_col126[5] <= 1'b0;
                    stage3_col126[6] <= 1'b0;
                    stage3_col126[7] <= 1'b0;
                    stage3_col126[8] <= 1'b0;
                    stage3_col126[9] <= 1'b0;
                    stage3_col126[10] <= 1'b0;
                    stage3_col127[0] <= 1'b0;
                    stage3_col127[1] <= 1'b0;
                    stage3_col127[2] <= 1'b0;
                    stage3_col127[3] <= 1'b0;
                    stage3_col127[4] <= 1'b0;
                    stage3_col127[5] <= 1'b0;
                    stage3_col127[6] <= 1'b0;
                    stage3_col127[7] <= 1'b0;
                    stage3_col127[8] <= 1'b0;
                    stage3_col127[9] <= 1'b0;
                    stage3_col127[10] <= 1'b0;
                    stage3_col127[11] <= 1'b0;
                    stage3_col127[12] <= 1'b0;
                    stage3_col127[13] <= 1'b0;
                    stage3_col127[14] <= 1'b0;
                    stage3_col127[15] <= 1'b0;
                    stage3_col127[16] <= 1'b0;
                    stage3_col127[17] <= 1'b0;
                    stage3_col127[18] <= 1'b0;
                    stage3_col127[19] <= 1'b0;
                    stage3_col127[20] <= 1'b0;
                    stage3_col127[21] <= 1'b0;
                    stage3_col127[22] <= 1'b0;
                    stage3_col127[23] <= 1'b0;
                    stage3_col127[24] <= 1'b0;
                    stage3_col127[25] <= 1'b0;
                    stage3_col127[26] <= 1'b0;
                    stage3_col127[27] <= 1'b0;
                    stage3_col127[28] <= 1'b0;
                    stage3_col127[29] <= 1'b0;
                    stage3_col127[30] <= 1'b0;
                    stage3_col127[31] <= 1'b0;
                    stage3_col127[32] <= 1'b0;
                    stage3_col127[33] <= 1'b0;
                    stage3_col127[34] <= 1'b0;
                    stage3_col127[35] <= 1'b0;
                    stage3_col127[36] <= 1'b0;
                    stage3_col127[37] <= 1'b0;
                    stage3_col127[38] <= 1'b0;
                    stage3_col127[39] <= 1'b0;
                    stage3_col127[40] <= 1'b0;
                    stage3_col127[41] <= 1'b0;
                    stage3_col127[42] <= 1'b0;
                    stage3_col127[43] <= 1'b0;
                    stage3_col127[44] <= 1'b0;
                    stage3_col127[45] <= 1'b0;
                    stage3_col127[46] <= 1'b0;
                    stage3_col127[47] <= 1'b0;
                    stage3_col127[48] <= 1'b0;
                    stage3_col127[49] <= 1'b0;
                    stage3_col127[50] <= 1'b0;
                    stage3_col127[51] <= 1'b0;
                    stage3_col127[52] <= 1'b0;
                    stage3_col127[53] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage3_col0[0] <= stage2_col0[0];
                    stage3_col1[0] <= stage2_col1[0];
                    stage3_col2[0] <= ha_s2_c2_n0_s;
                    stage3_col3[0] <= ha_s2_c2_n0_c;
                    stage3_col3[1] <= stage2_col3[0];
                    stage3_col4[0] <= fa_s2_c4_n0_s;
                    stage3_col5[0] <= fa_s2_c4_n0_c;
                    stage3_col5[1] <= stage2_col5[0];
                    stage3_col5[2] <= stage2_col5[1];
                    stage3_col6[0] <= stage2_col6[0];
                    stage3_col6[1] <= stage2_col6[1];
                    stage3_col7[0] <= stage2_col7[0];
                    stage3_col7[1] <= stage2_col7[1];
                    stage3_col8[0] <= stage2_col8[0];
                    stage3_col8[1] <= stage2_col8[1];
                    stage3_col9[0] <= fa_s2_c9_n1_s;
                    stage3_col9[1] <= stage2_col9[3];
                    stage3_col10[0] <= fa_s2_c9_n1_c;
                    stage3_col10[1] <= fa_s2_c10_n2_s;
                    stage3_col11[0] <= fa_s2_c10_n2_c;
                    stage3_col11[1] <= fa_s2_c11_n3_s;
                    stage3_col12[0] <= fa_s2_c11_n3_c;
                    stage3_col12[1] <= fa_s2_c12_n4_s;
                    stage3_col13[0] <= fa_s2_c12_n4_c;
                    stage3_col13[1] <= fa_s2_c13_n5_s;
                    stage3_col13[2] <= stage2_col13[3];
                    stage3_col13[3] <= stage2_col13[4];
                    stage3_col14[0] <= fa_s2_c13_n5_c;
                    stage3_col14[1] <= fa_s2_c14_n6_s;
                    stage3_col14[2] <= stage2_col14[3];
                    stage3_col15[0] <= fa_s2_c14_n6_c;
                    stage3_col15[1] <= fa_s2_c15_n7_s;
                    stage3_col15[2] <= stage2_col15[3];
                    stage3_col16[0] <= fa_s2_c15_n7_c;
                    stage3_col16[1] <= fa_s2_c16_n8_s;
                    stage3_col16[2] <= stage2_col16[3];
                    stage3_col17[0] <= fa_s2_c16_n8_c;
                    stage3_col17[1] <= fa_s2_c17_n9_s;
                    stage3_col17[2] <= stage2_col17[3];
                    stage3_col18[0] <= fa_s2_c17_n9_c;
                    stage3_col18[1] <= fa_s2_c18_n10_s;
                    stage3_col18[2] <= fa_s2_c18_n11_s;
                    stage3_col19[0] <= fa_s2_c18_n10_c;
                    stage3_col19[1] <= fa_s2_c18_n11_c;
                    stage3_col19[2] <= fa_s2_c19_n12_s;
                    stage3_col19[3] <= stage2_col19[3];
                    stage3_col19[4] <= stage2_col19[4];
                    stage3_col20[0] <= fa_s2_c19_n12_c;
                    stage3_col20[1] <= fa_s2_c20_n13_s;
                    stage3_col20[2] <= stage2_col20[3];
                    stage3_col20[3] <= stage2_col20[4];
                    stage3_col21[0] <= fa_s2_c20_n13_c;
                    stage3_col21[1] <= fa_s2_c21_n14_s;
                    stage3_col21[2] <= stage2_col21[3];
                    stage3_col21[3] <= stage2_col21[4];
                    stage3_col22[0] <= fa_s2_c21_n14_c;
                    stage3_col22[1] <= fa_s2_c22_n15_s;
                    stage3_col22[2] <= fa_s2_c22_n16_s;
                    stage3_col22[3] <= stage2_col22[6];
                    stage3_col23[0] <= fa_s2_c22_n15_c;
                    stage3_col23[1] <= fa_s2_c22_n16_c;
                    stage3_col23[2] <= fa_s2_c23_n17_s;
                    stage3_col23[3] <= fa_s2_c23_n18_s;
                    stage3_col24[0] <= fa_s2_c23_n17_c;
                    stage3_col24[1] <= fa_s2_c23_n18_c;
                    stage3_col24[2] <= fa_s2_c24_n19_s;
                    stage3_col24[3] <= fa_s2_c24_n20_s;
                    stage3_col25[0] <= fa_s2_c24_n19_c;
                    stage3_col25[1] <= fa_s2_c24_n20_c;
                    stage3_col25[2] <= fa_s2_c25_n21_s;
                    stage3_col25[3] <= fa_s2_c25_n22_s;
                    stage3_col26[0] <= fa_s2_c25_n21_c;
                    stage3_col26[1] <= fa_s2_c25_n22_c;
                    stage3_col26[2] <= fa_s2_c26_n23_s;
                    stage3_col26[3] <= fa_s2_c26_n24_s;
                    stage3_col27[0] <= fa_s2_c26_n23_c;
                    stage3_col27[1] <= fa_s2_c26_n24_c;
                    stage3_col27[2] <= fa_s2_c27_n25_s;
                    stage3_col27[3] <= fa_s2_c27_n26_s;
                    stage3_col27[4] <= stage2_col27[6];
                    stage3_col27[5] <= stage2_col27[7];
                    stage3_col28[0] <= fa_s2_c27_n25_c;
                    stage3_col28[1] <= fa_s2_c27_n26_c;
                    stage3_col28[2] <= fa_s2_c28_n27_s;
                    stage3_col28[3] <= fa_s2_c28_n28_s;
                    stage3_col28[4] <= stage2_col28[6];
                    stage3_col29[0] <= fa_s2_c28_n27_c;
                    stage3_col29[1] <= fa_s2_c28_n28_c;
                    stage3_col29[2] <= fa_s2_c29_n29_s;
                    stage3_col29[3] <= fa_s2_c29_n30_s;
                    stage3_col29[4] <= stage2_col29[6];
                    stage3_col30[0] <= fa_s2_c29_n29_c;
                    stage3_col30[1] <= fa_s2_c29_n30_c;
                    stage3_col30[2] <= fa_s2_c30_n31_s;
                    stage3_col30[3] <= fa_s2_c30_n32_s;
                    stage3_col30[4] <= stage2_col30[6];
                    stage3_col31[0] <= fa_s2_c30_n31_c;
                    stage3_col31[1] <= fa_s2_c30_n32_c;
                    stage3_col31[2] <= fa_s2_c31_n33_s;
                    stage3_col31[3] <= fa_s2_c31_n34_s;
                    stage3_col31[4] <= fa_s2_c31_n35_s;
                    stage3_col32[0] <= fa_s2_c31_n33_c;
                    stage3_col32[1] <= fa_s2_c31_n34_c;
                    stage3_col32[2] <= fa_s2_c31_n35_c;
                    stage3_col32[3] <= fa_s2_c32_n36_s;
                    stage3_col32[4] <= fa_s2_c32_n37_s;
                    stage3_col32[5] <= stage2_col32[6];
                    stage3_col32[6] <= stage2_col32[7];
                    stage3_col33[0] <= fa_s2_c32_n36_c;
                    stage3_col33[1] <= fa_s2_c32_n37_c;
                    stage3_col33[2] <= fa_s2_c33_n38_s;
                    stage3_col33[3] <= fa_s2_c33_n39_s;
                    stage3_col33[4] <= stage2_col33[6];
                    stage3_col33[5] <= stage2_col33[7];
                    stage3_col34[0] <= fa_s2_c33_n38_c;
                    stage3_col34[1] <= fa_s2_c33_n39_c;
                    stage3_col34[2] <= fa_s2_c34_n40_s;
                    stage3_col34[3] <= fa_s2_c34_n41_s;
                    stage3_col34[4] <= stage2_col34[6];
                    stage3_col34[5] <= stage2_col34[7];
                    stage3_col35[0] <= fa_s2_c34_n40_c;
                    stage3_col35[1] <= fa_s2_c34_n41_c;
                    stage3_col35[2] <= fa_s2_c35_n42_s;
                    stage3_col35[3] <= fa_s2_c35_n43_s;
                    stage3_col35[4] <= stage2_col35[6];
                    stage3_col35[5] <= stage2_col35[7];
                    stage3_col36[0] <= fa_s2_c35_n42_c;
                    stage3_col36[1] <= fa_s2_c35_n43_c;
                    stage3_col36[2] <= fa_s2_c36_n44_s;
                    stage3_col36[3] <= fa_s2_c36_n45_s;
                    stage3_col36[4] <= fa_s2_c36_n46_s;
                    stage3_col36[5] <= stage2_col36[9];
                    stage3_col37[0] <= fa_s2_c36_n44_c;
                    stage3_col37[1] <= fa_s2_c36_n45_c;
                    stage3_col37[2] <= fa_s2_c36_n46_c;
                    stage3_col37[3] <= fa_s2_c37_n47_s;
                    stage3_col37[4] <= fa_s2_c37_n48_s;
                    stage3_col37[5] <= fa_s2_c37_n49_s;
                    stage3_col38[0] <= fa_s2_c37_n47_c;
                    stage3_col38[1] <= fa_s2_c37_n48_c;
                    stage3_col38[2] <= fa_s2_c37_n49_c;
                    stage3_col38[3] <= fa_s2_c38_n50_s;
                    stage3_col38[4] <= fa_s2_c38_n51_s;
                    stage3_col38[5] <= fa_s2_c38_n52_s;
                    stage3_col39[0] <= fa_s2_c38_n50_c;
                    stage3_col39[1] <= fa_s2_c38_n51_c;
                    stage3_col39[2] <= fa_s2_c38_n52_c;
                    stage3_col39[3] <= fa_s2_c39_n53_s;
                    stage3_col39[4] <= fa_s2_c39_n54_s;
                    stage3_col39[5] <= fa_s2_c39_n55_s;
                    stage3_col40[0] <= fa_s2_c39_n53_c;
                    stage3_col40[1] <= fa_s2_c39_n54_c;
                    stage3_col40[2] <= fa_s2_c39_n55_c;
                    stage3_col40[3] <= fa_s2_c40_n56_s;
                    stage3_col40[4] <= fa_s2_c40_n57_s;
                    stage3_col40[5] <= fa_s2_c40_n58_s;
                    stage3_col40[6] <= stage2_col40[9];
                    stage3_col40[7] <= stage2_col40[10];
                    stage3_col41[0] <= fa_s2_c40_n56_c;
                    stage3_col41[1] <= fa_s2_c40_n57_c;
                    stage3_col41[2] <= fa_s2_c40_n58_c;
                    stage3_col41[3] <= fa_s2_c41_n59_s;
                    stage3_col41[4] <= fa_s2_c41_n60_s;
                    stage3_col41[5] <= fa_s2_c41_n61_s;
                    stage3_col41[6] <= stage2_col41[9];
                    stage3_col42[0] <= fa_s2_c41_n59_c;
                    stage3_col42[1] <= fa_s2_c41_n60_c;
                    stage3_col42[2] <= fa_s2_c41_n61_c;
                    stage3_col42[3] <= fa_s2_c42_n62_s;
                    stage3_col42[4] <= fa_s2_c42_n63_s;
                    stage3_col42[5] <= fa_s2_c42_n64_s;
                    stage3_col42[6] <= stage2_col42[9];
                    stage3_col43[0] <= fa_s2_c42_n62_c;
                    stage3_col43[1] <= fa_s2_c42_n63_c;
                    stage3_col43[2] <= fa_s2_c42_n64_c;
                    stage3_col43[3] <= fa_s2_c43_n65_s;
                    stage3_col43[4] <= fa_s2_c43_n66_s;
                    stage3_col43[5] <= fa_s2_c43_n67_s;
                    stage3_col43[6] <= stage2_col43[9];
                    stage3_col44[0] <= fa_s2_c43_n65_c;
                    stage3_col44[1] <= fa_s2_c43_n66_c;
                    stage3_col44[2] <= fa_s2_c43_n67_c;
                    stage3_col44[3] <= fa_s2_c44_n68_s;
                    stage3_col44[4] <= fa_s2_c44_n69_s;
                    stage3_col44[5] <= fa_s2_c44_n70_s;
                    stage3_col44[6] <= stage2_col44[9];
                    stage3_col45[0] <= fa_s2_c44_n68_c;
                    stage3_col45[1] <= fa_s2_c44_n69_c;
                    stage3_col45[2] <= fa_s2_c44_n70_c;
                    stage3_col45[3] <= fa_s2_c45_n71_s;
                    stage3_col45[4] <= fa_s2_c45_n72_s;
                    stage3_col45[5] <= fa_s2_c45_n73_s;
                    stage3_col45[6] <= fa_s2_c45_n74_s;
                    stage3_col46[0] <= fa_s2_c45_n71_c;
                    stage3_col46[1] <= fa_s2_c45_n72_c;
                    stage3_col46[2] <= fa_s2_c45_n73_c;
                    stage3_col46[3] <= fa_s2_c45_n74_c;
                    stage3_col46[4] <= fa_s2_c46_n75_s;
                    stage3_col46[5] <= fa_s2_c46_n76_s;
                    stage3_col46[6] <= fa_s2_c46_n77_s;
                    stage3_col46[7] <= stage2_col46[9];
                    stage3_col46[8] <= stage2_col46[10];
                    stage3_col47[0] <= fa_s2_c46_n75_c;
                    stage3_col47[1] <= fa_s2_c46_n76_c;
                    stage3_col47[2] <= fa_s2_c46_n77_c;
                    stage3_col47[3] <= fa_s2_c47_n78_s;
                    stage3_col47[4] <= fa_s2_c47_n79_s;
                    stage3_col47[5] <= fa_s2_c47_n80_s;
                    stage3_col47[6] <= stage2_col47[9];
                    stage3_col47[7] <= stage2_col47[10];
                    stage3_col48[0] <= fa_s2_c47_n78_c;
                    stage3_col48[1] <= fa_s2_c47_n79_c;
                    stage3_col48[2] <= fa_s2_c47_n80_c;
                    stage3_col48[3] <= fa_s2_c48_n81_s;
                    stage3_col48[4] <= fa_s2_c48_n82_s;
                    stage3_col48[5] <= fa_s2_c48_n83_s;
                    stage3_col48[6] <= stage2_col48[9];
                    stage3_col48[7] <= stage2_col48[10];
                    stage3_col49[0] <= fa_s2_c48_n81_c;
                    stage3_col49[1] <= fa_s2_c48_n82_c;
                    stage3_col49[2] <= fa_s2_c48_n83_c;
                    stage3_col49[3] <= fa_s2_c49_n84_s;
                    stage3_col49[4] <= fa_s2_c49_n85_s;
                    stage3_col49[5] <= fa_s2_c49_n86_s;
                    stage3_col49[6] <= fa_s2_c49_n87_s;
                    stage3_col49[7] <= stage2_col49[12];
                    stage3_col50[0] <= fa_s2_c49_n84_c;
                    stage3_col50[1] <= fa_s2_c49_n85_c;
                    stage3_col50[2] <= fa_s2_c49_n86_c;
                    stage3_col50[3] <= fa_s2_c49_n87_c;
                    stage3_col50[4] <= fa_s2_c50_n88_s;
                    stage3_col50[5] <= fa_s2_c50_n89_s;
                    stage3_col50[6] <= fa_s2_c50_n90_s;
                    stage3_col50[7] <= fa_s2_c50_n91_s;
                    stage3_col51[0] <= fa_s2_c50_n88_c;
                    stage3_col51[1] <= fa_s2_c50_n89_c;
                    stage3_col51[2] <= fa_s2_c50_n90_c;
                    stage3_col51[3] <= fa_s2_c50_n91_c;
                    stage3_col51[4] <= fa_s2_c51_n92_s;
                    stage3_col51[5] <= fa_s2_c51_n93_s;
                    stage3_col51[6] <= fa_s2_c51_n94_s;
                    stage3_col51[7] <= fa_s2_c51_n95_s;
                    stage3_col52[0] <= fa_s2_c51_n92_c;
                    stage3_col52[1] <= fa_s2_c51_n93_c;
                    stage3_col52[2] <= fa_s2_c51_n94_c;
                    stage3_col52[3] <= fa_s2_c51_n95_c;
                    stage3_col52[4] <= fa_s2_c52_n96_s;
                    stage3_col52[5] <= fa_s2_c52_n97_s;
                    stage3_col52[6] <= fa_s2_c52_n98_s;
                    stage3_col52[7] <= fa_s2_c52_n99_s;
                    stage3_col53[0] <= fa_s2_c52_n96_c;
                    stage3_col53[1] <= fa_s2_c52_n97_c;
                    stage3_col53[2] <= fa_s2_c52_n98_c;
                    stage3_col53[3] <= fa_s2_c52_n99_c;
                    stage3_col53[4] <= fa_s2_c53_n100_s;
                    stage3_col53[5] <= fa_s2_c53_n101_s;
                    stage3_col53[6] <= fa_s2_c53_n102_s;
                    stage3_col53[7] <= fa_s2_c53_n103_s;
                    stage3_col54[0] <= fa_s2_c53_n100_c;
                    stage3_col54[1] <= fa_s2_c53_n101_c;
                    stage3_col54[2] <= fa_s2_c53_n102_c;
                    stage3_col54[3] <= fa_s2_c53_n103_c;
                    stage3_col54[4] <= fa_s2_c54_n104_s;
                    stage3_col54[5] <= fa_s2_c54_n105_s;
                    stage3_col54[6] <= fa_s2_c54_n106_s;
                    stage3_col54[7] <= fa_s2_c54_n107_s;
                    stage3_col54[8] <= stage2_col54[12];
                    stage3_col54[9] <= stage2_col54[13];
                    stage3_col55[0] <= fa_s2_c54_n104_c;
                    stage3_col55[1] <= fa_s2_c54_n105_c;
                    stage3_col55[2] <= fa_s2_c54_n106_c;
                    stage3_col55[3] <= fa_s2_c54_n107_c;
                    stage3_col55[4] <= fa_s2_c55_n108_s;
                    stage3_col55[5] <= fa_s2_c55_n109_s;
                    stage3_col55[6] <= fa_s2_c55_n110_s;
                    stage3_col55[7] <= fa_s2_c55_n111_s;
                    stage3_col55[8] <= stage2_col55[12];
                    stage3_col56[0] <= fa_s2_c55_n108_c;
                    stage3_col56[1] <= fa_s2_c55_n109_c;
                    stage3_col56[2] <= fa_s2_c55_n110_c;
                    stage3_col56[3] <= fa_s2_c55_n111_c;
                    stage3_col56[4] <= fa_s2_c56_n112_s;
                    stage3_col56[5] <= fa_s2_c56_n113_s;
                    stage3_col56[6] <= fa_s2_c56_n114_s;
                    stage3_col56[7] <= fa_s2_c56_n115_s;
                    stage3_col56[8] <= stage2_col56[12];
                    stage3_col57[0] <= fa_s2_c56_n112_c;
                    stage3_col57[1] <= fa_s2_c56_n113_c;
                    stage3_col57[2] <= fa_s2_c56_n114_c;
                    stage3_col57[3] <= fa_s2_c56_n115_c;
                    stage3_col57[4] <= fa_s2_c57_n116_s;
                    stage3_col57[5] <= fa_s2_c57_n117_s;
                    stage3_col57[6] <= fa_s2_c57_n118_s;
                    stage3_col57[7] <= fa_s2_c57_n119_s;
                    stage3_col57[8] <= stage2_col57[12];
                    stage3_col58[0] <= fa_s2_c57_n116_c;
                    stage3_col58[1] <= fa_s2_c57_n117_c;
                    stage3_col58[2] <= fa_s2_c57_n118_c;
                    stage3_col58[3] <= fa_s2_c57_n119_c;
                    stage3_col58[4] <= fa_s2_c58_n120_s;
                    stage3_col58[5] <= fa_s2_c58_n121_s;
                    stage3_col58[6] <= fa_s2_c58_n122_s;
                    stage3_col58[7] <= fa_s2_c58_n123_s;
                    stage3_col58[8] <= fa_s2_c58_n124_s;
                    stage3_col59[0] <= fa_s2_c58_n120_c;
                    stage3_col59[1] <= fa_s2_c58_n121_c;
                    stage3_col59[2] <= fa_s2_c58_n122_c;
                    stage3_col59[3] <= fa_s2_c58_n123_c;
                    stage3_col59[4] <= fa_s2_c58_n124_c;
                    stage3_col59[5] <= fa_s2_c59_n125_s;
                    stage3_col59[6] <= fa_s2_c59_n126_s;
                    stage3_col59[7] <= fa_s2_c59_n127_s;
                    stage3_col59[8] <= fa_s2_c59_n128_s;
                    stage3_col59[9] <= stage2_col59[12];
                    stage3_col59[10] <= stage2_col59[13];
                    stage3_col60[0] <= fa_s2_c59_n125_c;
                    stage3_col60[1] <= fa_s2_c59_n126_c;
                    stage3_col60[2] <= fa_s2_c59_n127_c;
                    stage3_col60[3] <= fa_s2_c59_n128_c;
                    stage3_col60[4] <= fa_s2_c60_n129_s;
                    stage3_col60[5] <= fa_s2_c60_n130_s;
                    stage3_col60[6] <= fa_s2_c60_n131_s;
                    stage3_col60[7] <= fa_s2_c60_n132_s;
                    stage3_col60[8] <= stage2_col60[12];
                    stage3_col60[9] <= stage2_col60[13];
                    stage3_col61[0] <= fa_s2_c60_n129_c;
                    stage3_col61[1] <= fa_s2_c60_n130_c;
                    stage3_col61[2] <= fa_s2_c60_n131_c;
                    stage3_col61[3] <= fa_s2_c60_n132_c;
                    stage3_col61[4] <= fa_s2_c61_n133_s;
                    stage3_col61[5] <= fa_s2_c61_n134_s;
                    stage3_col61[6] <= fa_s2_c61_n135_s;
                    stage3_col61[7] <= fa_s2_c61_n136_s;
                    stage3_col61[8] <= stage2_col61[12];
                    stage3_col61[9] <= stage2_col61[13];
                    stage3_col62[0] <= fa_s2_c61_n133_c;
                    stage3_col62[1] <= fa_s2_c61_n134_c;
                    stage3_col62[2] <= fa_s2_c61_n135_c;
                    stage3_col62[3] <= fa_s2_c61_n136_c;
                    stage3_col62[4] <= fa_s2_c62_n137_s;
                    stage3_col62[5] <= fa_s2_c62_n138_s;
                    stage3_col62[6] <= fa_s2_c62_n139_s;
                    stage3_col62[7] <= fa_s2_c62_n140_s;
                    stage3_col62[8] <= stage2_col62[12];
                    stage3_col62[9] <= stage2_col62[13];
                    stage3_col63[0] <= fa_s2_c62_n137_c;
                    stage3_col63[1] <= fa_s2_c62_n138_c;
                    stage3_col63[2] <= fa_s2_c62_n139_c;
                    stage3_col63[3] <= fa_s2_c62_n140_c;
                    stage3_col63[4] <= fa_s2_c63_n141_s;
                    stage3_col63[5] <= fa_s2_c63_n142_s;
                    stage3_col63[6] <= fa_s2_c63_n143_s;
                    stage3_col63[7] <= fa_s2_c63_n144_s;
                    stage3_col63[8] <= fa_s2_c63_n145_s;
                    stage3_col63[9] <= stage2_col63[15];
                    stage3_col64[0] <= fa_s2_c63_n141_c;
                    stage3_col64[1] <= fa_s2_c63_n142_c;
                    stage3_col64[2] <= fa_s2_c63_n143_c;
                    stage3_col64[3] <= fa_s2_c63_n144_c;
                    stage3_col64[4] <= fa_s2_c63_n145_c;
                    stage3_col64[5] <= fa_s2_c64_n146_s;
                    stage3_col64[6] <= fa_s2_c64_n147_s;
                    stage3_col64[7] <= fa_s2_c64_n148_s;
                    stage3_col64[8] <= fa_s2_c64_n149_s;
                    stage3_col64[9] <= stage2_col64[12];
                    stage3_col64[10] <= stage2_col64[13];
                    stage3_col65[0] <= fa_s2_c64_n146_c;
                    stage3_col65[1] <= fa_s2_c64_n147_c;
                    stage3_col65[2] <= fa_s2_c64_n148_c;
                    stage3_col65[3] <= fa_s2_c64_n149_c;
                    stage3_col65[4] <= fa_s2_c65_n150_s;
                    stage3_col65[5] <= fa_s2_c65_n151_s;
                    stage3_col65[6] <= fa_s2_c65_n152_s;
                    stage3_col65[7] <= fa_s2_c65_n153_s;
                    stage3_col65[8] <= fa_s2_c65_n154_s;
                    stage3_col65[9] <= stage2_col65[15];
                    stage3_col66[0] <= fa_s2_c65_n150_c;
                    stage3_col66[1] <= fa_s2_c65_n151_c;
                    stage3_col66[2] <= fa_s2_c65_n152_c;
                    stage3_col66[3] <= fa_s2_c65_n153_c;
                    stage3_col66[4] <= fa_s2_c65_n154_c;
                    stage3_col66[5] <= fa_s2_c66_n155_s;
                    stage3_col66[6] <= fa_s2_c66_n156_s;
                    stage3_col66[7] <= fa_s2_c66_n157_s;
                    stage3_col66[8] <= fa_s2_c66_n158_s;
                    stage3_col66[9] <= stage2_col66[12];
                    stage3_col66[10] <= stage2_col66[13];
                    stage3_col67[0] <= fa_s2_c66_n155_c;
                    stage3_col67[1] <= fa_s2_c66_n156_c;
                    stage3_col67[2] <= fa_s2_c66_n157_c;
                    stage3_col67[3] <= fa_s2_c66_n158_c;
                    stage3_col67[4] <= fa_s2_c67_n159_s;
                    stage3_col67[5] <= fa_s2_c67_n160_s;
                    stage3_col67[6] <= fa_s2_c67_n161_s;
                    stage3_col67[7] <= fa_s2_c67_n162_s;
                    stage3_col67[8] <= fa_s2_c67_n163_s;
                    stage3_col67[9] <= stage2_col67[15];
                    stage3_col68[0] <= fa_s2_c67_n159_c;
                    stage3_col68[1] <= fa_s2_c67_n160_c;
                    stage3_col68[2] <= fa_s2_c67_n161_c;
                    stage3_col68[3] <= fa_s2_c67_n162_c;
                    stage3_col68[4] <= fa_s2_c67_n163_c;
                    stage3_col68[5] <= fa_s2_c68_n164_s;
                    stage3_col68[6] <= fa_s2_c68_n165_s;
                    stage3_col68[7] <= fa_s2_c68_n166_s;
                    stage3_col68[8] <= fa_s2_c68_n167_s;
                    stage3_col68[9] <= stage2_col68[12];
                    stage3_col68[10] <= stage2_col68[13];
                    stage3_col69[0] <= fa_s2_c68_n164_c;
                    stage3_col69[1] <= fa_s2_c68_n165_c;
                    stage3_col69[2] <= fa_s2_c68_n166_c;
                    stage3_col69[3] <= fa_s2_c68_n167_c;
                    stage3_col69[4] <= fa_s2_c69_n168_s;
                    stage3_col69[5] <= fa_s2_c69_n169_s;
                    stage3_col69[6] <= fa_s2_c69_n170_s;
                    stage3_col69[7] <= fa_s2_c69_n171_s;
                    stage3_col69[8] <= fa_s2_c69_n172_s;
                    stage3_col69[9] <= stage2_col69[15];
                    stage3_col70[0] <= fa_s2_c69_n168_c;
                    stage3_col70[1] <= fa_s2_c69_n169_c;
                    stage3_col70[2] <= fa_s2_c69_n170_c;
                    stage3_col70[3] <= fa_s2_c69_n171_c;
                    stage3_col70[4] <= fa_s2_c69_n172_c;
                    stage3_col70[5] <= fa_s2_c70_n173_s;
                    stage3_col70[6] <= fa_s2_c70_n174_s;
                    stage3_col70[7] <= fa_s2_c70_n175_s;
                    stage3_col70[8] <= fa_s2_c70_n176_s;
                    stage3_col70[9] <= stage2_col70[12];
                    stage3_col70[10] <= stage2_col70[13];
                    stage3_col71[0] <= fa_s2_c70_n173_c;
                    stage3_col71[1] <= fa_s2_c70_n174_c;
                    stage3_col71[2] <= fa_s2_c70_n175_c;
                    stage3_col71[3] <= fa_s2_c70_n176_c;
                    stage3_col71[4] <= fa_s2_c71_n177_s;
                    stage3_col71[5] <= fa_s2_c71_n178_s;
                    stage3_col71[6] <= fa_s2_c71_n179_s;
                    stage3_col71[7] <= fa_s2_c71_n180_s;
                    stage3_col71[8] <= fa_s2_c71_n181_s;
                    stage3_col71[9] <= stage2_col71[15];
                    stage3_col72[0] <= fa_s2_c71_n177_c;
                    stage3_col72[1] <= fa_s2_c71_n178_c;
                    stage3_col72[2] <= fa_s2_c71_n179_c;
                    stage3_col72[3] <= fa_s2_c71_n180_c;
                    stage3_col72[4] <= fa_s2_c71_n181_c;
                    stage3_col72[5] <= fa_s2_c72_n182_s;
                    stage3_col72[6] <= fa_s2_c72_n183_s;
                    stage3_col72[7] <= fa_s2_c72_n184_s;
                    stage3_col72[8] <= fa_s2_c72_n185_s;
                    stage3_col72[9] <= stage2_col72[12];
                    stage3_col72[10] <= stage2_col72[13];
                    stage3_col73[0] <= fa_s2_c72_n182_c;
                    stage3_col73[1] <= fa_s2_c72_n183_c;
                    stage3_col73[2] <= fa_s2_c72_n184_c;
                    stage3_col73[3] <= fa_s2_c72_n185_c;
                    stage3_col73[4] <= fa_s2_c73_n186_s;
                    stage3_col73[5] <= fa_s2_c73_n187_s;
                    stage3_col73[6] <= fa_s2_c73_n188_s;
                    stage3_col73[7] <= fa_s2_c73_n189_s;
                    stage3_col73[8] <= fa_s2_c73_n190_s;
                    stage3_col73[9] <= stage2_col73[15];
                    stage3_col74[0] <= fa_s2_c73_n186_c;
                    stage3_col74[1] <= fa_s2_c73_n187_c;
                    stage3_col74[2] <= fa_s2_c73_n188_c;
                    stage3_col74[3] <= fa_s2_c73_n189_c;
                    stage3_col74[4] <= fa_s2_c73_n190_c;
                    stage3_col74[5] <= fa_s2_c74_n191_s;
                    stage3_col74[6] <= fa_s2_c74_n192_s;
                    stage3_col74[7] <= fa_s2_c74_n193_s;
                    stage3_col74[8] <= fa_s2_c74_n194_s;
                    stage3_col74[9] <= stage2_col74[12];
                    stage3_col74[10] <= stage2_col74[13];
                    stage3_col75[0] <= fa_s2_c74_n191_c;
                    stage3_col75[1] <= fa_s2_c74_n192_c;
                    stage3_col75[2] <= fa_s2_c74_n193_c;
                    stage3_col75[3] <= fa_s2_c74_n194_c;
                    stage3_col75[4] <= fa_s2_c75_n195_s;
                    stage3_col75[5] <= fa_s2_c75_n196_s;
                    stage3_col75[6] <= fa_s2_c75_n197_s;
                    stage3_col75[7] <= fa_s2_c75_n198_s;
                    stage3_col75[8] <= fa_s2_c75_n199_s;
                    stage3_col75[9] <= stage2_col75[15];
                    stage3_col76[0] <= fa_s2_c75_n195_c;
                    stage3_col76[1] <= fa_s2_c75_n196_c;
                    stage3_col76[2] <= fa_s2_c75_n197_c;
                    stage3_col76[3] <= fa_s2_c75_n198_c;
                    stage3_col76[4] <= fa_s2_c75_n199_c;
                    stage3_col76[5] <= fa_s2_c76_n200_s;
                    stage3_col76[6] <= fa_s2_c76_n201_s;
                    stage3_col76[7] <= fa_s2_c76_n202_s;
                    stage3_col76[8] <= fa_s2_c76_n203_s;
                    stage3_col76[9] <= stage2_col76[12];
                    stage3_col76[10] <= stage2_col76[13];
                    stage3_col77[0] <= fa_s2_c76_n200_c;
                    stage3_col77[1] <= fa_s2_c76_n201_c;
                    stage3_col77[2] <= fa_s2_c76_n202_c;
                    stage3_col77[3] <= fa_s2_c76_n203_c;
                    stage3_col77[4] <= fa_s2_c77_n204_s;
                    stage3_col77[5] <= fa_s2_c77_n205_s;
                    stage3_col77[6] <= fa_s2_c77_n206_s;
                    stage3_col77[7] <= fa_s2_c77_n207_s;
                    stage3_col77[8] <= fa_s2_c77_n208_s;
                    stage3_col77[9] <= stage2_col77[15];
                    stage3_col78[0] <= fa_s2_c77_n204_c;
                    stage3_col78[1] <= fa_s2_c77_n205_c;
                    stage3_col78[2] <= fa_s2_c77_n206_c;
                    stage3_col78[3] <= fa_s2_c77_n207_c;
                    stage3_col78[4] <= fa_s2_c77_n208_c;
                    stage3_col78[5] <= fa_s2_c78_n209_s;
                    stage3_col78[6] <= fa_s2_c78_n210_s;
                    stage3_col78[7] <= fa_s2_c78_n211_s;
                    stage3_col78[8] <= fa_s2_c78_n212_s;
                    stage3_col78[9] <= stage2_col78[12];
                    stage3_col78[10] <= stage2_col78[13];
                    stage3_col79[0] <= fa_s2_c78_n209_c;
                    stage3_col79[1] <= fa_s2_c78_n210_c;
                    stage3_col79[2] <= fa_s2_c78_n211_c;
                    stage3_col79[3] <= fa_s2_c78_n212_c;
                    stage3_col79[4] <= fa_s2_c79_n213_s;
                    stage3_col79[5] <= fa_s2_c79_n214_s;
                    stage3_col79[6] <= fa_s2_c79_n215_s;
                    stage3_col79[7] <= fa_s2_c79_n216_s;
                    stage3_col79[8] <= fa_s2_c79_n217_s;
                    stage3_col79[9] <= stage2_col79[15];
                    stage3_col80[0] <= fa_s2_c79_n213_c;
                    stage3_col80[1] <= fa_s2_c79_n214_c;
                    stage3_col80[2] <= fa_s2_c79_n215_c;
                    stage3_col80[3] <= fa_s2_c79_n216_c;
                    stage3_col80[4] <= fa_s2_c79_n217_c;
                    stage3_col80[5] <= fa_s2_c80_n218_s;
                    stage3_col80[6] <= fa_s2_c80_n219_s;
                    stage3_col80[7] <= fa_s2_c80_n220_s;
                    stage3_col80[8] <= fa_s2_c80_n221_s;
                    stage3_col80[9] <= stage2_col80[12];
                    stage3_col80[10] <= stage2_col80[13];
                    stage3_col81[0] <= fa_s2_c80_n218_c;
                    stage3_col81[1] <= fa_s2_c80_n219_c;
                    stage3_col81[2] <= fa_s2_c80_n220_c;
                    stage3_col81[3] <= fa_s2_c80_n221_c;
                    stage3_col81[4] <= fa_s2_c81_n222_s;
                    stage3_col81[5] <= fa_s2_c81_n223_s;
                    stage3_col81[6] <= fa_s2_c81_n224_s;
                    stage3_col81[7] <= fa_s2_c81_n225_s;
                    stage3_col81[8] <= fa_s2_c81_n226_s;
                    stage3_col81[9] <= stage2_col81[15];
                    stage3_col82[0] <= fa_s2_c81_n222_c;
                    stage3_col82[1] <= fa_s2_c81_n223_c;
                    stage3_col82[2] <= fa_s2_c81_n224_c;
                    stage3_col82[3] <= fa_s2_c81_n225_c;
                    stage3_col82[4] <= fa_s2_c81_n226_c;
                    stage3_col82[5] <= fa_s2_c82_n227_s;
                    stage3_col82[6] <= fa_s2_c82_n228_s;
                    stage3_col82[7] <= fa_s2_c82_n229_s;
                    stage3_col82[8] <= fa_s2_c82_n230_s;
                    stage3_col82[9] <= stage2_col82[12];
                    stage3_col82[10] <= stage2_col82[13];
                    stage3_col83[0] <= fa_s2_c82_n227_c;
                    stage3_col83[1] <= fa_s2_c82_n228_c;
                    stage3_col83[2] <= fa_s2_c82_n229_c;
                    stage3_col83[3] <= fa_s2_c82_n230_c;
                    stage3_col83[4] <= fa_s2_c83_n231_s;
                    stage3_col83[5] <= fa_s2_c83_n232_s;
                    stage3_col83[6] <= fa_s2_c83_n233_s;
                    stage3_col83[7] <= fa_s2_c83_n234_s;
                    stage3_col83[8] <= fa_s2_c83_n235_s;
                    stage3_col83[9] <= stage2_col83[15];
                    stage3_col84[0] <= fa_s2_c83_n231_c;
                    stage3_col84[1] <= fa_s2_c83_n232_c;
                    stage3_col84[2] <= fa_s2_c83_n233_c;
                    stage3_col84[3] <= fa_s2_c83_n234_c;
                    stage3_col84[4] <= fa_s2_c83_n235_c;
                    stage3_col84[5] <= fa_s2_c84_n236_s;
                    stage3_col84[6] <= fa_s2_c84_n237_s;
                    stage3_col84[7] <= fa_s2_c84_n238_s;
                    stage3_col84[8] <= fa_s2_c84_n239_s;
                    stage3_col84[9] <= stage2_col84[12];
                    stage3_col84[10] <= stage2_col84[13];
                    stage3_col85[0] <= fa_s2_c84_n236_c;
                    stage3_col85[1] <= fa_s2_c84_n237_c;
                    stage3_col85[2] <= fa_s2_c84_n238_c;
                    stage3_col85[3] <= fa_s2_c84_n239_c;
                    stage3_col85[4] <= fa_s2_c85_n240_s;
                    stage3_col85[5] <= fa_s2_c85_n241_s;
                    stage3_col85[6] <= fa_s2_c85_n242_s;
                    stage3_col85[7] <= fa_s2_c85_n243_s;
                    stage3_col85[8] <= fa_s2_c85_n244_s;
                    stage3_col85[9] <= stage2_col85[15];
                    stage3_col86[0] <= fa_s2_c85_n240_c;
                    stage3_col86[1] <= fa_s2_c85_n241_c;
                    stage3_col86[2] <= fa_s2_c85_n242_c;
                    stage3_col86[3] <= fa_s2_c85_n243_c;
                    stage3_col86[4] <= fa_s2_c85_n244_c;
                    stage3_col86[5] <= fa_s2_c86_n245_s;
                    stage3_col86[6] <= fa_s2_c86_n246_s;
                    stage3_col86[7] <= fa_s2_c86_n247_s;
                    stage3_col86[8] <= fa_s2_c86_n248_s;
                    stage3_col86[9] <= stage2_col86[12];
                    stage3_col86[10] <= stage2_col86[13];
                    stage3_col87[0] <= fa_s2_c86_n245_c;
                    stage3_col87[1] <= fa_s2_c86_n246_c;
                    stage3_col87[2] <= fa_s2_c86_n247_c;
                    stage3_col87[3] <= fa_s2_c86_n248_c;
                    stage3_col87[4] <= fa_s2_c87_n249_s;
                    stage3_col87[5] <= fa_s2_c87_n250_s;
                    stage3_col87[6] <= fa_s2_c87_n251_s;
                    stage3_col87[7] <= fa_s2_c87_n252_s;
                    stage3_col87[8] <= fa_s2_c87_n253_s;
                    stage3_col87[9] <= stage2_col87[15];
                    stage3_col88[0] <= fa_s2_c87_n249_c;
                    stage3_col88[1] <= fa_s2_c87_n250_c;
                    stage3_col88[2] <= fa_s2_c87_n251_c;
                    stage3_col88[3] <= fa_s2_c87_n252_c;
                    stage3_col88[4] <= fa_s2_c87_n253_c;
                    stage3_col88[5] <= fa_s2_c88_n254_s;
                    stage3_col88[6] <= fa_s2_c88_n255_s;
                    stage3_col88[7] <= fa_s2_c88_n256_s;
                    stage3_col88[8] <= fa_s2_c88_n257_s;
                    stage3_col88[9] <= stage2_col88[12];
                    stage3_col88[10] <= stage2_col88[13];
                    stage3_col89[0] <= fa_s2_c88_n254_c;
                    stage3_col89[1] <= fa_s2_c88_n255_c;
                    stage3_col89[2] <= fa_s2_c88_n256_c;
                    stage3_col89[3] <= fa_s2_c88_n257_c;
                    stage3_col89[4] <= fa_s2_c89_n258_s;
                    stage3_col89[5] <= fa_s2_c89_n259_s;
                    stage3_col89[6] <= fa_s2_c89_n260_s;
                    stage3_col89[7] <= fa_s2_c89_n261_s;
                    stage3_col89[8] <= fa_s2_c89_n262_s;
                    stage3_col89[9] <= stage2_col89[15];
                    stage3_col90[0] <= fa_s2_c89_n258_c;
                    stage3_col90[1] <= fa_s2_c89_n259_c;
                    stage3_col90[2] <= fa_s2_c89_n260_c;
                    stage3_col90[3] <= fa_s2_c89_n261_c;
                    stage3_col90[4] <= fa_s2_c89_n262_c;
                    stage3_col90[5] <= fa_s2_c90_n263_s;
                    stage3_col90[6] <= fa_s2_c90_n264_s;
                    stage3_col90[7] <= fa_s2_c90_n265_s;
                    stage3_col90[8] <= fa_s2_c90_n266_s;
                    stage3_col90[9] <= stage2_col90[12];
                    stage3_col90[10] <= stage2_col90[13];
                    stage3_col91[0] <= fa_s2_c90_n263_c;
                    stage3_col91[1] <= fa_s2_c90_n264_c;
                    stage3_col91[2] <= fa_s2_c90_n265_c;
                    stage3_col91[3] <= fa_s2_c90_n266_c;
                    stage3_col91[4] <= fa_s2_c91_n267_s;
                    stage3_col91[5] <= fa_s2_c91_n268_s;
                    stage3_col91[6] <= fa_s2_c91_n269_s;
                    stage3_col91[7] <= fa_s2_c91_n270_s;
                    stage3_col91[8] <= fa_s2_c91_n271_s;
                    stage3_col91[9] <= stage2_col91[15];
                    stage3_col92[0] <= fa_s2_c91_n267_c;
                    stage3_col92[1] <= fa_s2_c91_n268_c;
                    stage3_col92[2] <= fa_s2_c91_n269_c;
                    stage3_col92[3] <= fa_s2_c91_n270_c;
                    stage3_col92[4] <= fa_s2_c91_n271_c;
                    stage3_col92[5] <= fa_s2_c92_n272_s;
                    stage3_col92[6] <= fa_s2_c92_n273_s;
                    stage3_col92[7] <= fa_s2_c92_n274_s;
                    stage3_col92[8] <= fa_s2_c92_n275_s;
                    stage3_col92[9] <= stage2_col92[12];
                    stage3_col92[10] <= stage2_col92[13];
                    stage3_col93[0] <= fa_s2_c92_n272_c;
                    stage3_col93[1] <= fa_s2_c92_n273_c;
                    stage3_col93[2] <= fa_s2_c92_n274_c;
                    stage3_col93[3] <= fa_s2_c92_n275_c;
                    stage3_col93[4] <= fa_s2_c93_n276_s;
                    stage3_col93[5] <= fa_s2_c93_n277_s;
                    stage3_col93[6] <= fa_s2_c93_n278_s;
                    stage3_col93[7] <= fa_s2_c93_n279_s;
                    stage3_col93[8] <= fa_s2_c93_n280_s;
                    stage3_col93[9] <= stage2_col93[15];
                    stage3_col94[0] <= fa_s2_c93_n276_c;
                    stage3_col94[1] <= fa_s2_c93_n277_c;
                    stage3_col94[2] <= fa_s2_c93_n278_c;
                    stage3_col94[3] <= fa_s2_c93_n279_c;
                    stage3_col94[4] <= fa_s2_c93_n280_c;
                    stage3_col94[5] <= fa_s2_c94_n281_s;
                    stage3_col94[6] <= fa_s2_c94_n282_s;
                    stage3_col94[7] <= fa_s2_c94_n283_s;
                    stage3_col94[8] <= fa_s2_c94_n284_s;
                    stage3_col94[9] <= stage2_col94[12];
                    stage3_col94[10] <= stage2_col94[13];
                    stage3_col95[0] <= fa_s2_c94_n281_c;
                    stage3_col95[1] <= fa_s2_c94_n282_c;
                    stage3_col95[2] <= fa_s2_c94_n283_c;
                    stage3_col95[3] <= fa_s2_c94_n284_c;
                    stage3_col95[4] <= fa_s2_c95_n285_s;
                    stage3_col95[5] <= fa_s2_c95_n286_s;
                    stage3_col95[6] <= fa_s2_c95_n287_s;
                    stage3_col95[7] <= fa_s2_c95_n288_s;
                    stage3_col95[8] <= fa_s2_c95_n289_s;
                    stage3_col95[9] <= stage2_col95[15];
                    stage3_col96[0] <= fa_s2_c95_n285_c;
                    stage3_col96[1] <= fa_s2_c95_n286_c;
                    stage3_col96[2] <= fa_s2_c95_n287_c;
                    stage3_col96[3] <= fa_s2_c95_n288_c;
                    stage3_col96[4] <= fa_s2_c95_n289_c;
                    stage3_col96[5] <= fa_s2_c96_n290_s;
                    stage3_col96[6] <= fa_s2_c96_n291_s;
                    stage3_col96[7] <= fa_s2_c96_n292_s;
                    stage3_col96[8] <= fa_s2_c96_n293_s;
                    stage3_col96[9] <= stage2_col96[12];
                    stage3_col96[10] <= stage2_col96[13];
                    stage3_col97[0] <= fa_s2_c96_n290_c;
                    stage3_col97[1] <= fa_s2_c96_n291_c;
                    stage3_col97[2] <= fa_s2_c96_n292_c;
                    stage3_col97[3] <= fa_s2_c96_n293_c;
                    stage3_col97[4] <= fa_s2_c97_n294_s;
                    stage3_col97[5] <= fa_s2_c97_n295_s;
                    stage3_col97[6] <= fa_s2_c97_n296_s;
                    stage3_col97[7] <= fa_s2_c97_n297_s;
                    stage3_col97[8] <= fa_s2_c97_n298_s;
                    stage3_col97[9] <= stage2_col97[15];
                    stage3_col98[0] <= fa_s2_c97_n294_c;
                    stage3_col98[1] <= fa_s2_c97_n295_c;
                    stage3_col98[2] <= fa_s2_c97_n296_c;
                    stage3_col98[3] <= fa_s2_c97_n297_c;
                    stage3_col98[4] <= fa_s2_c97_n298_c;
                    stage3_col98[5] <= fa_s2_c98_n299_s;
                    stage3_col98[6] <= fa_s2_c98_n300_s;
                    stage3_col98[7] <= fa_s2_c98_n301_s;
                    stage3_col98[8] <= fa_s2_c98_n302_s;
                    stage3_col98[9] <= stage2_col98[12];
                    stage3_col98[10] <= stage2_col98[13];
                    stage3_col99[0] <= fa_s2_c98_n299_c;
                    stage3_col99[1] <= fa_s2_c98_n300_c;
                    stage3_col99[2] <= fa_s2_c98_n301_c;
                    stage3_col99[3] <= fa_s2_c98_n302_c;
                    stage3_col99[4] <= fa_s2_c99_n303_s;
                    stage3_col99[5] <= fa_s2_c99_n304_s;
                    stage3_col99[6] <= fa_s2_c99_n305_s;
                    stage3_col99[7] <= fa_s2_c99_n306_s;
                    stage3_col99[8] <= fa_s2_c99_n307_s;
                    stage3_col99[9] <= stage2_col99[15];
                    stage3_col100[0] <= fa_s2_c99_n303_c;
                    stage3_col100[1] <= fa_s2_c99_n304_c;
                    stage3_col100[2] <= fa_s2_c99_n305_c;
                    stage3_col100[3] <= fa_s2_c99_n306_c;
                    stage3_col100[4] <= fa_s2_c99_n307_c;
                    stage3_col100[5] <= fa_s2_c100_n308_s;
                    stage3_col100[6] <= fa_s2_c100_n309_s;
                    stage3_col100[7] <= fa_s2_c100_n310_s;
                    stage3_col100[8] <= fa_s2_c100_n311_s;
                    stage3_col100[9] <= stage2_col100[12];
                    stage3_col100[10] <= stage2_col100[13];
                    stage3_col101[0] <= fa_s2_c100_n308_c;
                    stage3_col101[1] <= fa_s2_c100_n309_c;
                    stage3_col101[2] <= fa_s2_c100_n310_c;
                    stage3_col101[3] <= fa_s2_c100_n311_c;
                    stage3_col101[4] <= fa_s2_c101_n312_s;
                    stage3_col101[5] <= fa_s2_c101_n313_s;
                    stage3_col101[6] <= fa_s2_c101_n314_s;
                    stage3_col101[7] <= fa_s2_c101_n315_s;
                    stage3_col101[8] <= fa_s2_c101_n316_s;
                    stage3_col101[9] <= stage2_col101[15];
                    stage3_col102[0] <= fa_s2_c101_n312_c;
                    stage3_col102[1] <= fa_s2_c101_n313_c;
                    stage3_col102[2] <= fa_s2_c101_n314_c;
                    stage3_col102[3] <= fa_s2_c101_n315_c;
                    stage3_col102[4] <= fa_s2_c101_n316_c;
                    stage3_col102[5] <= fa_s2_c102_n317_s;
                    stage3_col102[6] <= fa_s2_c102_n318_s;
                    stage3_col102[7] <= fa_s2_c102_n319_s;
                    stage3_col102[8] <= fa_s2_c102_n320_s;
                    stage3_col102[9] <= stage2_col102[12];
                    stage3_col102[10] <= stage2_col102[13];
                    stage3_col103[0] <= fa_s2_c102_n317_c;
                    stage3_col103[1] <= fa_s2_c102_n318_c;
                    stage3_col103[2] <= fa_s2_c102_n319_c;
                    stage3_col103[3] <= fa_s2_c102_n320_c;
                    stage3_col103[4] <= fa_s2_c103_n321_s;
                    stage3_col103[5] <= fa_s2_c103_n322_s;
                    stage3_col103[6] <= fa_s2_c103_n323_s;
                    stage3_col103[7] <= fa_s2_c103_n324_s;
                    stage3_col103[8] <= fa_s2_c103_n325_s;
                    stage3_col103[9] <= stage2_col103[15];
                    stage3_col104[0] <= fa_s2_c103_n321_c;
                    stage3_col104[1] <= fa_s2_c103_n322_c;
                    stage3_col104[2] <= fa_s2_c103_n323_c;
                    stage3_col104[3] <= fa_s2_c103_n324_c;
                    stage3_col104[4] <= fa_s2_c103_n325_c;
                    stage3_col104[5] <= fa_s2_c104_n326_s;
                    stage3_col104[6] <= fa_s2_c104_n327_s;
                    stage3_col104[7] <= fa_s2_c104_n328_s;
                    stage3_col104[8] <= fa_s2_c104_n329_s;
                    stage3_col104[9] <= stage2_col104[12];
                    stage3_col104[10] <= stage2_col104[13];
                    stage3_col105[0] <= fa_s2_c104_n326_c;
                    stage3_col105[1] <= fa_s2_c104_n327_c;
                    stage3_col105[2] <= fa_s2_c104_n328_c;
                    stage3_col105[3] <= fa_s2_c104_n329_c;
                    stage3_col105[4] <= fa_s2_c105_n330_s;
                    stage3_col105[5] <= fa_s2_c105_n331_s;
                    stage3_col105[6] <= fa_s2_c105_n332_s;
                    stage3_col105[7] <= fa_s2_c105_n333_s;
                    stage3_col105[8] <= fa_s2_c105_n334_s;
                    stage3_col105[9] <= stage2_col105[15];
                    stage3_col106[0] <= fa_s2_c105_n330_c;
                    stage3_col106[1] <= fa_s2_c105_n331_c;
                    stage3_col106[2] <= fa_s2_c105_n332_c;
                    stage3_col106[3] <= fa_s2_c105_n333_c;
                    stage3_col106[4] <= fa_s2_c105_n334_c;
                    stage3_col106[5] <= fa_s2_c106_n335_s;
                    stage3_col106[6] <= fa_s2_c106_n336_s;
                    stage3_col106[7] <= fa_s2_c106_n337_s;
                    stage3_col106[8] <= fa_s2_c106_n338_s;
                    stage3_col106[9] <= stage2_col106[12];
                    stage3_col106[10] <= stage2_col106[13];
                    stage3_col107[0] <= fa_s2_c106_n335_c;
                    stage3_col107[1] <= fa_s2_c106_n336_c;
                    stage3_col107[2] <= fa_s2_c106_n337_c;
                    stage3_col107[3] <= fa_s2_c106_n338_c;
                    stage3_col107[4] <= fa_s2_c107_n339_s;
                    stage3_col107[5] <= fa_s2_c107_n340_s;
                    stage3_col107[6] <= fa_s2_c107_n341_s;
                    stage3_col107[7] <= fa_s2_c107_n342_s;
                    stage3_col107[8] <= fa_s2_c107_n343_s;
                    stage3_col107[9] <= stage2_col107[15];
                    stage3_col108[0] <= fa_s2_c107_n339_c;
                    stage3_col108[1] <= fa_s2_c107_n340_c;
                    stage3_col108[2] <= fa_s2_c107_n341_c;
                    stage3_col108[3] <= fa_s2_c107_n342_c;
                    stage3_col108[4] <= fa_s2_c107_n343_c;
                    stage3_col108[5] <= fa_s2_c108_n344_s;
                    stage3_col108[6] <= fa_s2_c108_n345_s;
                    stage3_col108[7] <= fa_s2_c108_n346_s;
                    stage3_col108[8] <= fa_s2_c108_n347_s;
                    stage3_col108[9] <= stage2_col108[12];
                    stage3_col108[10] <= stage2_col108[13];
                    stage3_col109[0] <= fa_s2_c108_n344_c;
                    stage3_col109[1] <= fa_s2_c108_n345_c;
                    stage3_col109[2] <= fa_s2_c108_n346_c;
                    stage3_col109[3] <= fa_s2_c108_n347_c;
                    stage3_col109[4] <= fa_s2_c109_n348_s;
                    stage3_col109[5] <= fa_s2_c109_n349_s;
                    stage3_col109[6] <= fa_s2_c109_n350_s;
                    stage3_col109[7] <= fa_s2_c109_n351_s;
                    stage3_col109[8] <= fa_s2_c109_n352_s;
                    stage3_col109[9] <= stage2_col109[15];
                    stage3_col110[0] <= fa_s2_c109_n348_c;
                    stage3_col110[1] <= fa_s2_c109_n349_c;
                    stage3_col110[2] <= fa_s2_c109_n350_c;
                    stage3_col110[3] <= fa_s2_c109_n351_c;
                    stage3_col110[4] <= fa_s2_c109_n352_c;
                    stage3_col110[5] <= fa_s2_c110_n353_s;
                    stage3_col110[6] <= fa_s2_c110_n354_s;
                    stage3_col110[7] <= fa_s2_c110_n355_s;
                    stage3_col110[8] <= fa_s2_c110_n356_s;
                    stage3_col110[9] <= stage2_col110[12];
                    stage3_col110[10] <= stage2_col110[13];
                    stage3_col111[0] <= fa_s2_c110_n353_c;
                    stage3_col111[1] <= fa_s2_c110_n354_c;
                    stage3_col111[2] <= fa_s2_c110_n355_c;
                    stage3_col111[3] <= fa_s2_c110_n356_c;
                    stage3_col111[4] <= fa_s2_c111_n357_s;
                    stage3_col111[5] <= fa_s2_c111_n358_s;
                    stage3_col111[6] <= fa_s2_c111_n359_s;
                    stage3_col111[7] <= fa_s2_c111_n360_s;
                    stage3_col111[8] <= fa_s2_c111_n361_s;
                    stage3_col111[9] <= stage2_col111[15];
                    stage3_col112[0] <= fa_s2_c111_n357_c;
                    stage3_col112[1] <= fa_s2_c111_n358_c;
                    stage3_col112[2] <= fa_s2_c111_n359_c;
                    stage3_col112[3] <= fa_s2_c111_n360_c;
                    stage3_col112[4] <= fa_s2_c111_n361_c;
                    stage3_col112[5] <= fa_s2_c112_n362_s;
                    stage3_col112[6] <= fa_s2_c112_n363_s;
                    stage3_col112[7] <= fa_s2_c112_n364_s;
                    stage3_col112[8] <= fa_s2_c112_n365_s;
                    stage3_col112[9] <= stage2_col112[12];
                    stage3_col112[10] <= stage2_col112[13];
                    stage3_col113[0] <= fa_s2_c112_n362_c;
                    stage3_col113[1] <= fa_s2_c112_n363_c;
                    stage3_col113[2] <= fa_s2_c112_n364_c;
                    stage3_col113[3] <= fa_s2_c112_n365_c;
                    stage3_col113[4] <= fa_s2_c113_n366_s;
                    stage3_col113[5] <= fa_s2_c113_n367_s;
                    stage3_col113[6] <= fa_s2_c113_n368_s;
                    stage3_col113[7] <= fa_s2_c113_n369_s;
                    stage3_col113[8] <= fa_s2_c113_n370_s;
                    stage3_col113[9] <= stage2_col113[15];
                    stage3_col114[0] <= fa_s2_c113_n366_c;
                    stage3_col114[1] <= fa_s2_c113_n367_c;
                    stage3_col114[2] <= fa_s2_c113_n368_c;
                    stage3_col114[3] <= fa_s2_c113_n369_c;
                    stage3_col114[4] <= fa_s2_c113_n370_c;
                    stage3_col114[5] <= fa_s2_c114_n371_s;
                    stage3_col114[6] <= fa_s2_c114_n372_s;
                    stage3_col114[7] <= fa_s2_c114_n373_s;
                    stage3_col114[8] <= fa_s2_c114_n374_s;
                    stage3_col114[9] <= stage2_col114[12];
                    stage3_col114[10] <= stage2_col114[13];
                    stage3_col115[0] <= fa_s2_c114_n371_c;
                    stage3_col115[1] <= fa_s2_c114_n372_c;
                    stage3_col115[2] <= fa_s2_c114_n373_c;
                    stage3_col115[3] <= fa_s2_c114_n374_c;
                    stage3_col115[4] <= fa_s2_c115_n375_s;
                    stage3_col115[5] <= fa_s2_c115_n376_s;
                    stage3_col115[6] <= fa_s2_c115_n377_s;
                    stage3_col115[7] <= fa_s2_c115_n378_s;
                    stage3_col115[8] <= fa_s2_c115_n379_s;
                    stage3_col115[9] <= stage2_col115[15];
                    stage3_col116[0] <= fa_s2_c115_n375_c;
                    stage3_col116[1] <= fa_s2_c115_n376_c;
                    stage3_col116[2] <= fa_s2_c115_n377_c;
                    stage3_col116[3] <= fa_s2_c115_n378_c;
                    stage3_col116[4] <= fa_s2_c115_n379_c;
                    stage3_col116[5] <= fa_s2_c116_n380_s;
                    stage3_col116[6] <= fa_s2_c116_n381_s;
                    stage3_col116[7] <= fa_s2_c116_n382_s;
                    stage3_col116[8] <= fa_s2_c116_n383_s;
                    stage3_col116[9] <= stage2_col116[12];
                    stage3_col116[10] <= stage2_col116[13];
                    stage3_col117[0] <= fa_s2_c116_n380_c;
                    stage3_col117[1] <= fa_s2_c116_n381_c;
                    stage3_col117[2] <= fa_s2_c116_n382_c;
                    stage3_col117[3] <= fa_s2_c116_n383_c;
                    stage3_col117[4] <= fa_s2_c117_n384_s;
                    stage3_col117[5] <= fa_s2_c117_n385_s;
                    stage3_col117[6] <= fa_s2_c117_n386_s;
                    stage3_col117[7] <= fa_s2_c117_n387_s;
                    stage3_col117[8] <= fa_s2_c117_n388_s;
                    stage3_col117[9] <= stage2_col117[15];
                    stage3_col118[0] <= fa_s2_c117_n384_c;
                    stage3_col118[1] <= fa_s2_c117_n385_c;
                    stage3_col118[2] <= fa_s2_c117_n386_c;
                    stage3_col118[3] <= fa_s2_c117_n387_c;
                    stage3_col118[4] <= fa_s2_c117_n388_c;
                    stage3_col118[5] <= fa_s2_c118_n389_s;
                    stage3_col118[6] <= fa_s2_c118_n390_s;
                    stage3_col118[7] <= fa_s2_c118_n391_s;
                    stage3_col118[8] <= fa_s2_c118_n392_s;
                    stage3_col118[9] <= stage2_col118[12];
                    stage3_col118[10] <= stage2_col118[13];
                    stage3_col119[0] <= fa_s2_c118_n389_c;
                    stage3_col119[1] <= fa_s2_c118_n390_c;
                    stage3_col119[2] <= fa_s2_c118_n391_c;
                    stage3_col119[3] <= fa_s2_c118_n392_c;
                    stage3_col119[4] <= fa_s2_c119_n393_s;
                    stage3_col119[5] <= fa_s2_c119_n394_s;
                    stage3_col119[6] <= fa_s2_c119_n395_s;
                    stage3_col119[7] <= fa_s2_c119_n396_s;
                    stage3_col119[8] <= fa_s2_c119_n397_s;
                    stage3_col119[9] <= stage2_col119[15];
                    stage3_col120[0] <= fa_s2_c119_n393_c;
                    stage3_col120[1] <= fa_s2_c119_n394_c;
                    stage3_col120[2] <= fa_s2_c119_n395_c;
                    stage3_col120[3] <= fa_s2_c119_n396_c;
                    stage3_col120[4] <= fa_s2_c119_n397_c;
                    stage3_col120[5] <= fa_s2_c120_n398_s;
                    stage3_col120[6] <= fa_s2_c120_n399_s;
                    stage3_col120[7] <= fa_s2_c120_n400_s;
                    stage3_col120[8] <= fa_s2_c120_n401_s;
                    stage3_col120[9] <= stage2_col120[12];
                    stage3_col120[10] <= stage2_col120[13];
                    stage3_col121[0] <= fa_s2_c120_n398_c;
                    stage3_col121[1] <= fa_s2_c120_n399_c;
                    stage3_col121[2] <= fa_s2_c120_n400_c;
                    stage3_col121[3] <= fa_s2_c120_n401_c;
                    stage3_col121[4] <= fa_s2_c121_n402_s;
                    stage3_col121[5] <= fa_s2_c121_n403_s;
                    stage3_col121[6] <= fa_s2_c121_n404_s;
                    stage3_col121[7] <= fa_s2_c121_n405_s;
                    stage3_col121[8] <= fa_s2_c121_n406_s;
                    stage3_col121[9] <= stage2_col121[15];
                    stage3_col122[0] <= fa_s2_c121_n402_c;
                    stage3_col122[1] <= fa_s2_c121_n403_c;
                    stage3_col122[2] <= fa_s2_c121_n404_c;
                    stage3_col122[3] <= fa_s2_c121_n405_c;
                    stage3_col122[4] <= fa_s2_c121_n406_c;
                    stage3_col122[5] <= fa_s2_c122_n407_s;
                    stage3_col122[6] <= fa_s2_c122_n408_s;
                    stage3_col122[7] <= fa_s2_c122_n409_s;
                    stage3_col122[8] <= fa_s2_c122_n410_s;
                    stage3_col122[9] <= stage2_col122[12];
                    stage3_col122[10] <= stage2_col122[13];
                    stage3_col123[0] <= fa_s2_c122_n407_c;
                    stage3_col123[1] <= fa_s2_c122_n408_c;
                    stage3_col123[2] <= fa_s2_c122_n409_c;
                    stage3_col123[3] <= fa_s2_c122_n410_c;
                    stage3_col123[4] <= fa_s2_c123_n411_s;
                    stage3_col123[5] <= fa_s2_c123_n412_s;
                    stage3_col123[6] <= fa_s2_c123_n413_s;
                    stage3_col123[7] <= fa_s2_c123_n414_s;
                    stage3_col123[8] <= fa_s2_c123_n415_s;
                    stage3_col123[9] <= stage2_col123[15];
                    stage3_col124[0] <= fa_s2_c123_n411_c;
                    stage3_col124[1] <= fa_s2_c123_n412_c;
                    stage3_col124[2] <= fa_s2_c123_n413_c;
                    stage3_col124[3] <= fa_s2_c123_n414_c;
                    stage3_col124[4] <= fa_s2_c123_n415_c;
                    stage3_col124[5] <= fa_s2_c124_n416_s;
                    stage3_col124[6] <= fa_s2_c124_n417_s;
                    stage3_col124[7] <= fa_s2_c124_n418_s;
                    stage3_col124[8] <= fa_s2_c124_n419_s;
                    stage3_col124[9] <= stage2_col124[12];
                    stage3_col124[10] <= stage2_col124[13];
                    stage3_col125[0] <= fa_s2_c124_n416_c;
                    stage3_col125[1] <= fa_s2_c124_n417_c;
                    stage3_col125[2] <= fa_s2_c124_n418_c;
                    stage3_col125[3] <= fa_s2_c124_n419_c;
                    stage3_col125[4] <= fa_s2_c125_n420_s;
                    stage3_col125[5] <= fa_s2_c125_n421_s;
                    stage3_col125[6] <= fa_s2_c125_n422_s;
                    stage3_col125[7] <= fa_s2_c125_n423_s;
                    stage3_col125[8] <= fa_s2_c125_n424_s;
                    stage3_col125[9] <= stage2_col125[15];
                    stage3_col126[0] <= fa_s2_c125_n420_c;
                    stage3_col126[1] <= fa_s2_c125_n421_c;
                    stage3_col126[2] <= fa_s2_c125_n422_c;
                    stage3_col126[3] <= fa_s2_c125_n423_c;
                    stage3_col126[4] <= fa_s2_c125_n424_c;
                    stage3_col126[5] <= fa_s2_c126_n425_s;
                    stage3_col126[6] <= fa_s2_c126_n426_s;
                    stage3_col126[7] <= fa_s2_c126_n427_s;
                    stage3_col126[8] <= fa_s2_c126_n428_s;
                    stage3_col126[9] <= stage2_col126[12];
                    stage3_col126[10] <= stage2_col126[13];
                    stage3_col127[0] <= fa_s2_c126_n425_c;
                    stage3_col127[1] <= fa_s2_c126_n426_c;
                    stage3_col127[2] <= fa_s2_c126_n427_c;
                    stage3_col127[3] <= fa_s2_c126_n428_c;
                    stage3_col127[4] <= stage2_col127[0];
                    stage3_col127[5] <= stage2_col127[1];
                    stage3_col127[6] <= stage2_col127[2];
                    stage3_col127[7] <= stage2_col127[3];
                    stage3_col127[8] <= stage2_col127[4];
                    stage3_col127[9] <= stage2_col127[5];
                    stage3_col127[10] <= stage2_col127[6];
                    stage3_col127[11] <= stage2_col127[7];
                    stage3_col127[12] <= stage2_col127[8];
                    stage3_col127[13] <= stage2_col127[9];
                    stage3_col127[14] <= stage2_col127[10];
                    stage3_col127[15] <= stage2_col127[11];
                    stage3_col127[16] <= stage2_col127[12];
                    stage3_col127[17] <= stage2_col127[13];
                    stage3_col127[18] <= stage2_col127[14];
                    stage3_col127[19] <= stage2_col127[15];
                    stage3_col127[20] <= stage2_col127[16];
                    stage3_col127[21] <= stage2_col127[17];
                    stage3_col127[22] <= stage2_col127[18];
                    stage3_col127[23] <= stage2_col127[18];
                    stage3_col127[24] <= stage2_col127[18];
                    stage3_col127[25] <= stage2_col127[18];
                    stage3_col127[26] <= stage2_col127[18];
                    stage3_col127[27] <= stage2_col127[18];
                    stage3_col127[28] <= stage2_col127[18];
                    stage3_col127[29] <= stage2_col127[18];
                    stage3_col127[30] <= stage2_col127[18];
                    stage3_col127[31] <= stage2_col127[18];
                    stage3_col127[32] <= stage2_col127[18];
                    stage3_col127[33] <= stage2_col127[18];
                    stage3_col127[34] <= stage2_col127[18];
                    stage3_col127[35] <= stage2_col127[18];
                    stage3_col127[36] <= stage2_col127[18];
                    stage3_col127[37] <= stage2_col127[18];
                    stage3_col127[38] <= stage2_col127[18];
                    stage3_col127[39] <= stage2_col127[18];
                    stage3_col127[40] <= stage2_col127[18];
                    stage3_col127[41] <= stage2_col127[18];
                    stage3_col127[42] <= stage2_col127[18];
                    stage3_col127[43] <= stage2_col127[18];
                    stage3_col127[44] <= stage2_col127[18];
                    stage3_col127[45] <= stage2_col127[18];
                    stage3_col127[46] <= stage2_col127[18];
                    stage3_col127[47] <= stage2_col127[18];
                    stage3_col127[48] <= stage2_col127[18];
                    stage3_col127[49] <= stage2_col127[18];
                    stage3_col127[50] <= stage2_col127[18];
                    stage3_col127[51] <= stage2_col127[18];
                    stage3_col127[52] <= stage2_col127[18];
                    stage3_col127[53] <= stage2_col127[18];
                end
            end
        end else begin : gen_stage3_no_pipe
            // Combinational assignment
            always_comb begin
                stage3_col0[0] = stage2_col0[0];
                stage3_col1[0] = stage2_col1[0];
                stage3_col2[0] = ha_s2_c2_n0_s;
                stage3_col3[0] = ha_s2_c2_n0_c;
                stage3_col3[1] = stage2_col3[0];
                stage3_col4[0] = fa_s2_c4_n0_s;
                stage3_col5[0] = fa_s2_c4_n0_c;
                stage3_col5[1] = stage2_col5[0];
                stage3_col5[2] = stage2_col5[1];
                stage3_col6[0] = stage2_col6[0];
                stage3_col6[1] = stage2_col6[1];
                stage3_col7[0] = stage2_col7[0];
                stage3_col7[1] = stage2_col7[1];
                stage3_col8[0] = stage2_col8[0];
                stage3_col8[1] = stage2_col8[1];
                stage3_col9[0] = fa_s2_c9_n1_s;
                stage3_col9[1] = stage2_col9[3];
                stage3_col10[0] = fa_s2_c9_n1_c;
                stage3_col10[1] = fa_s2_c10_n2_s;
                stage3_col11[0] = fa_s2_c10_n2_c;
                stage3_col11[1] = fa_s2_c11_n3_s;
                stage3_col12[0] = fa_s2_c11_n3_c;
                stage3_col12[1] = fa_s2_c12_n4_s;
                stage3_col13[0] = fa_s2_c12_n4_c;
                stage3_col13[1] = fa_s2_c13_n5_s;
                stage3_col13[2] = stage2_col13[3];
                stage3_col13[3] = stage2_col13[4];
                stage3_col14[0] = fa_s2_c13_n5_c;
                stage3_col14[1] = fa_s2_c14_n6_s;
                stage3_col14[2] = stage2_col14[3];
                stage3_col15[0] = fa_s2_c14_n6_c;
                stage3_col15[1] = fa_s2_c15_n7_s;
                stage3_col15[2] = stage2_col15[3];
                stage3_col16[0] = fa_s2_c15_n7_c;
                stage3_col16[1] = fa_s2_c16_n8_s;
                stage3_col16[2] = stage2_col16[3];
                stage3_col17[0] = fa_s2_c16_n8_c;
                stage3_col17[1] = fa_s2_c17_n9_s;
                stage3_col17[2] = stage2_col17[3];
                stage3_col18[0] = fa_s2_c17_n9_c;
                stage3_col18[1] = fa_s2_c18_n10_s;
                stage3_col18[2] = fa_s2_c18_n11_s;
                stage3_col19[0] = fa_s2_c18_n10_c;
                stage3_col19[1] = fa_s2_c18_n11_c;
                stage3_col19[2] = fa_s2_c19_n12_s;
                stage3_col19[3] = stage2_col19[3];
                stage3_col19[4] = stage2_col19[4];
                stage3_col20[0] = fa_s2_c19_n12_c;
                stage3_col20[1] = fa_s2_c20_n13_s;
                stage3_col20[2] = stage2_col20[3];
                stage3_col20[3] = stage2_col20[4];
                stage3_col21[0] = fa_s2_c20_n13_c;
                stage3_col21[1] = fa_s2_c21_n14_s;
                stage3_col21[2] = stage2_col21[3];
                stage3_col21[3] = stage2_col21[4];
                stage3_col22[0] = fa_s2_c21_n14_c;
                stage3_col22[1] = fa_s2_c22_n15_s;
                stage3_col22[2] = fa_s2_c22_n16_s;
                stage3_col22[3] = stage2_col22[6];
                stage3_col23[0] = fa_s2_c22_n15_c;
                stage3_col23[1] = fa_s2_c22_n16_c;
                stage3_col23[2] = fa_s2_c23_n17_s;
                stage3_col23[3] = fa_s2_c23_n18_s;
                stage3_col24[0] = fa_s2_c23_n17_c;
                stage3_col24[1] = fa_s2_c23_n18_c;
                stage3_col24[2] = fa_s2_c24_n19_s;
                stage3_col24[3] = fa_s2_c24_n20_s;
                stage3_col25[0] = fa_s2_c24_n19_c;
                stage3_col25[1] = fa_s2_c24_n20_c;
                stage3_col25[2] = fa_s2_c25_n21_s;
                stage3_col25[3] = fa_s2_c25_n22_s;
                stage3_col26[0] = fa_s2_c25_n21_c;
                stage3_col26[1] = fa_s2_c25_n22_c;
                stage3_col26[2] = fa_s2_c26_n23_s;
                stage3_col26[3] = fa_s2_c26_n24_s;
                stage3_col27[0] = fa_s2_c26_n23_c;
                stage3_col27[1] = fa_s2_c26_n24_c;
                stage3_col27[2] = fa_s2_c27_n25_s;
                stage3_col27[3] = fa_s2_c27_n26_s;
                stage3_col27[4] = stage2_col27[6];
                stage3_col27[5] = stage2_col27[7];
                stage3_col28[0] = fa_s2_c27_n25_c;
                stage3_col28[1] = fa_s2_c27_n26_c;
                stage3_col28[2] = fa_s2_c28_n27_s;
                stage3_col28[3] = fa_s2_c28_n28_s;
                stage3_col28[4] = stage2_col28[6];
                stage3_col29[0] = fa_s2_c28_n27_c;
                stage3_col29[1] = fa_s2_c28_n28_c;
                stage3_col29[2] = fa_s2_c29_n29_s;
                stage3_col29[3] = fa_s2_c29_n30_s;
                stage3_col29[4] = stage2_col29[6];
                stage3_col30[0] = fa_s2_c29_n29_c;
                stage3_col30[1] = fa_s2_c29_n30_c;
                stage3_col30[2] = fa_s2_c30_n31_s;
                stage3_col30[3] = fa_s2_c30_n32_s;
                stage3_col30[4] = stage2_col30[6];
                stage3_col31[0] = fa_s2_c30_n31_c;
                stage3_col31[1] = fa_s2_c30_n32_c;
                stage3_col31[2] = fa_s2_c31_n33_s;
                stage3_col31[3] = fa_s2_c31_n34_s;
                stage3_col31[4] = fa_s2_c31_n35_s;
                stage3_col32[0] = fa_s2_c31_n33_c;
                stage3_col32[1] = fa_s2_c31_n34_c;
                stage3_col32[2] = fa_s2_c31_n35_c;
                stage3_col32[3] = fa_s2_c32_n36_s;
                stage3_col32[4] = fa_s2_c32_n37_s;
                stage3_col32[5] = stage2_col32[6];
                stage3_col32[6] = stage2_col32[7];
                stage3_col33[0] = fa_s2_c32_n36_c;
                stage3_col33[1] = fa_s2_c32_n37_c;
                stage3_col33[2] = fa_s2_c33_n38_s;
                stage3_col33[3] = fa_s2_c33_n39_s;
                stage3_col33[4] = stage2_col33[6];
                stage3_col33[5] = stage2_col33[7];
                stage3_col34[0] = fa_s2_c33_n38_c;
                stage3_col34[1] = fa_s2_c33_n39_c;
                stage3_col34[2] = fa_s2_c34_n40_s;
                stage3_col34[3] = fa_s2_c34_n41_s;
                stage3_col34[4] = stage2_col34[6];
                stage3_col34[5] = stage2_col34[7];
                stage3_col35[0] = fa_s2_c34_n40_c;
                stage3_col35[1] = fa_s2_c34_n41_c;
                stage3_col35[2] = fa_s2_c35_n42_s;
                stage3_col35[3] = fa_s2_c35_n43_s;
                stage3_col35[4] = stage2_col35[6];
                stage3_col35[5] = stage2_col35[7];
                stage3_col36[0] = fa_s2_c35_n42_c;
                stage3_col36[1] = fa_s2_c35_n43_c;
                stage3_col36[2] = fa_s2_c36_n44_s;
                stage3_col36[3] = fa_s2_c36_n45_s;
                stage3_col36[4] = fa_s2_c36_n46_s;
                stage3_col36[5] = stage2_col36[9];
                stage3_col37[0] = fa_s2_c36_n44_c;
                stage3_col37[1] = fa_s2_c36_n45_c;
                stage3_col37[2] = fa_s2_c36_n46_c;
                stage3_col37[3] = fa_s2_c37_n47_s;
                stage3_col37[4] = fa_s2_c37_n48_s;
                stage3_col37[5] = fa_s2_c37_n49_s;
                stage3_col38[0] = fa_s2_c37_n47_c;
                stage3_col38[1] = fa_s2_c37_n48_c;
                stage3_col38[2] = fa_s2_c37_n49_c;
                stage3_col38[3] = fa_s2_c38_n50_s;
                stage3_col38[4] = fa_s2_c38_n51_s;
                stage3_col38[5] = fa_s2_c38_n52_s;
                stage3_col39[0] = fa_s2_c38_n50_c;
                stage3_col39[1] = fa_s2_c38_n51_c;
                stage3_col39[2] = fa_s2_c38_n52_c;
                stage3_col39[3] = fa_s2_c39_n53_s;
                stage3_col39[4] = fa_s2_c39_n54_s;
                stage3_col39[5] = fa_s2_c39_n55_s;
                stage3_col40[0] = fa_s2_c39_n53_c;
                stage3_col40[1] = fa_s2_c39_n54_c;
                stage3_col40[2] = fa_s2_c39_n55_c;
                stage3_col40[3] = fa_s2_c40_n56_s;
                stage3_col40[4] = fa_s2_c40_n57_s;
                stage3_col40[5] = fa_s2_c40_n58_s;
                stage3_col40[6] = stage2_col40[9];
                stage3_col40[7] = stage2_col40[10];
                stage3_col41[0] = fa_s2_c40_n56_c;
                stage3_col41[1] = fa_s2_c40_n57_c;
                stage3_col41[2] = fa_s2_c40_n58_c;
                stage3_col41[3] = fa_s2_c41_n59_s;
                stage3_col41[4] = fa_s2_c41_n60_s;
                stage3_col41[5] = fa_s2_c41_n61_s;
                stage3_col41[6] = stage2_col41[9];
                stage3_col42[0] = fa_s2_c41_n59_c;
                stage3_col42[1] = fa_s2_c41_n60_c;
                stage3_col42[2] = fa_s2_c41_n61_c;
                stage3_col42[3] = fa_s2_c42_n62_s;
                stage3_col42[4] = fa_s2_c42_n63_s;
                stage3_col42[5] = fa_s2_c42_n64_s;
                stage3_col42[6] = stage2_col42[9];
                stage3_col43[0] = fa_s2_c42_n62_c;
                stage3_col43[1] = fa_s2_c42_n63_c;
                stage3_col43[2] = fa_s2_c42_n64_c;
                stage3_col43[3] = fa_s2_c43_n65_s;
                stage3_col43[4] = fa_s2_c43_n66_s;
                stage3_col43[5] = fa_s2_c43_n67_s;
                stage3_col43[6] = stage2_col43[9];
                stage3_col44[0] = fa_s2_c43_n65_c;
                stage3_col44[1] = fa_s2_c43_n66_c;
                stage3_col44[2] = fa_s2_c43_n67_c;
                stage3_col44[3] = fa_s2_c44_n68_s;
                stage3_col44[4] = fa_s2_c44_n69_s;
                stage3_col44[5] = fa_s2_c44_n70_s;
                stage3_col44[6] = stage2_col44[9];
                stage3_col45[0] = fa_s2_c44_n68_c;
                stage3_col45[1] = fa_s2_c44_n69_c;
                stage3_col45[2] = fa_s2_c44_n70_c;
                stage3_col45[3] = fa_s2_c45_n71_s;
                stage3_col45[4] = fa_s2_c45_n72_s;
                stage3_col45[5] = fa_s2_c45_n73_s;
                stage3_col45[6] = fa_s2_c45_n74_s;
                stage3_col46[0] = fa_s2_c45_n71_c;
                stage3_col46[1] = fa_s2_c45_n72_c;
                stage3_col46[2] = fa_s2_c45_n73_c;
                stage3_col46[3] = fa_s2_c45_n74_c;
                stage3_col46[4] = fa_s2_c46_n75_s;
                stage3_col46[5] = fa_s2_c46_n76_s;
                stage3_col46[6] = fa_s2_c46_n77_s;
                stage3_col46[7] = stage2_col46[9];
                stage3_col46[8] = stage2_col46[10];
                stage3_col47[0] = fa_s2_c46_n75_c;
                stage3_col47[1] = fa_s2_c46_n76_c;
                stage3_col47[2] = fa_s2_c46_n77_c;
                stage3_col47[3] = fa_s2_c47_n78_s;
                stage3_col47[4] = fa_s2_c47_n79_s;
                stage3_col47[5] = fa_s2_c47_n80_s;
                stage3_col47[6] = stage2_col47[9];
                stage3_col47[7] = stage2_col47[10];
                stage3_col48[0] = fa_s2_c47_n78_c;
                stage3_col48[1] = fa_s2_c47_n79_c;
                stage3_col48[2] = fa_s2_c47_n80_c;
                stage3_col48[3] = fa_s2_c48_n81_s;
                stage3_col48[4] = fa_s2_c48_n82_s;
                stage3_col48[5] = fa_s2_c48_n83_s;
                stage3_col48[6] = stage2_col48[9];
                stage3_col48[7] = stage2_col48[10];
                stage3_col49[0] = fa_s2_c48_n81_c;
                stage3_col49[1] = fa_s2_c48_n82_c;
                stage3_col49[2] = fa_s2_c48_n83_c;
                stage3_col49[3] = fa_s2_c49_n84_s;
                stage3_col49[4] = fa_s2_c49_n85_s;
                stage3_col49[5] = fa_s2_c49_n86_s;
                stage3_col49[6] = fa_s2_c49_n87_s;
                stage3_col49[7] = stage2_col49[12];
                stage3_col50[0] = fa_s2_c49_n84_c;
                stage3_col50[1] = fa_s2_c49_n85_c;
                stage3_col50[2] = fa_s2_c49_n86_c;
                stage3_col50[3] = fa_s2_c49_n87_c;
                stage3_col50[4] = fa_s2_c50_n88_s;
                stage3_col50[5] = fa_s2_c50_n89_s;
                stage3_col50[6] = fa_s2_c50_n90_s;
                stage3_col50[7] = fa_s2_c50_n91_s;
                stage3_col51[0] = fa_s2_c50_n88_c;
                stage3_col51[1] = fa_s2_c50_n89_c;
                stage3_col51[2] = fa_s2_c50_n90_c;
                stage3_col51[3] = fa_s2_c50_n91_c;
                stage3_col51[4] = fa_s2_c51_n92_s;
                stage3_col51[5] = fa_s2_c51_n93_s;
                stage3_col51[6] = fa_s2_c51_n94_s;
                stage3_col51[7] = fa_s2_c51_n95_s;
                stage3_col52[0] = fa_s2_c51_n92_c;
                stage3_col52[1] = fa_s2_c51_n93_c;
                stage3_col52[2] = fa_s2_c51_n94_c;
                stage3_col52[3] = fa_s2_c51_n95_c;
                stage3_col52[4] = fa_s2_c52_n96_s;
                stage3_col52[5] = fa_s2_c52_n97_s;
                stage3_col52[6] = fa_s2_c52_n98_s;
                stage3_col52[7] = fa_s2_c52_n99_s;
                stage3_col53[0] = fa_s2_c52_n96_c;
                stage3_col53[1] = fa_s2_c52_n97_c;
                stage3_col53[2] = fa_s2_c52_n98_c;
                stage3_col53[3] = fa_s2_c52_n99_c;
                stage3_col53[4] = fa_s2_c53_n100_s;
                stage3_col53[5] = fa_s2_c53_n101_s;
                stage3_col53[6] = fa_s2_c53_n102_s;
                stage3_col53[7] = fa_s2_c53_n103_s;
                stage3_col54[0] = fa_s2_c53_n100_c;
                stage3_col54[1] = fa_s2_c53_n101_c;
                stage3_col54[2] = fa_s2_c53_n102_c;
                stage3_col54[3] = fa_s2_c53_n103_c;
                stage3_col54[4] = fa_s2_c54_n104_s;
                stage3_col54[5] = fa_s2_c54_n105_s;
                stage3_col54[6] = fa_s2_c54_n106_s;
                stage3_col54[7] = fa_s2_c54_n107_s;
                stage3_col54[8] = stage2_col54[12];
                stage3_col54[9] = stage2_col54[13];
                stage3_col55[0] = fa_s2_c54_n104_c;
                stage3_col55[1] = fa_s2_c54_n105_c;
                stage3_col55[2] = fa_s2_c54_n106_c;
                stage3_col55[3] = fa_s2_c54_n107_c;
                stage3_col55[4] = fa_s2_c55_n108_s;
                stage3_col55[5] = fa_s2_c55_n109_s;
                stage3_col55[6] = fa_s2_c55_n110_s;
                stage3_col55[7] = fa_s2_c55_n111_s;
                stage3_col55[8] = stage2_col55[12];
                stage3_col56[0] = fa_s2_c55_n108_c;
                stage3_col56[1] = fa_s2_c55_n109_c;
                stage3_col56[2] = fa_s2_c55_n110_c;
                stage3_col56[3] = fa_s2_c55_n111_c;
                stage3_col56[4] = fa_s2_c56_n112_s;
                stage3_col56[5] = fa_s2_c56_n113_s;
                stage3_col56[6] = fa_s2_c56_n114_s;
                stage3_col56[7] = fa_s2_c56_n115_s;
                stage3_col56[8] = stage2_col56[12];
                stage3_col57[0] = fa_s2_c56_n112_c;
                stage3_col57[1] = fa_s2_c56_n113_c;
                stage3_col57[2] = fa_s2_c56_n114_c;
                stage3_col57[3] = fa_s2_c56_n115_c;
                stage3_col57[4] = fa_s2_c57_n116_s;
                stage3_col57[5] = fa_s2_c57_n117_s;
                stage3_col57[6] = fa_s2_c57_n118_s;
                stage3_col57[7] = fa_s2_c57_n119_s;
                stage3_col57[8] = stage2_col57[12];
                stage3_col58[0] = fa_s2_c57_n116_c;
                stage3_col58[1] = fa_s2_c57_n117_c;
                stage3_col58[2] = fa_s2_c57_n118_c;
                stage3_col58[3] = fa_s2_c57_n119_c;
                stage3_col58[4] = fa_s2_c58_n120_s;
                stage3_col58[5] = fa_s2_c58_n121_s;
                stage3_col58[6] = fa_s2_c58_n122_s;
                stage3_col58[7] = fa_s2_c58_n123_s;
                stage3_col58[8] = fa_s2_c58_n124_s;
                stage3_col59[0] = fa_s2_c58_n120_c;
                stage3_col59[1] = fa_s2_c58_n121_c;
                stage3_col59[2] = fa_s2_c58_n122_c;
                stage3_col59[3] = fa_s2_c58_n123_c;
                stage3_col59[4] = fa_s2_c58_n124_c;
                stage3_col59[5] = fa_s2_c59_n125_s;
                stage3_col59[6] = fa_s2_c59_n126_s;
                stage3_col59[7] = fa_s2_c59_n127_s;
                stage3_col59[8] = fa_s2_c59_n128_s;
                stage3_col59[9] = stage2_col59[12];
                stage3_col59[10] = stage2_col59[13];
                stage3_col60[0] = fa_s2_c59_n125_c;
                stage3_col60[1] = fa_s2_c59_n126_c;
                stage3_col60[2] = fa_s2_c59_n127_c;
                stage3_col60[3] = fa_s2_c59_n128_c;
                stage3_col60[4] = fa_s2_c60_n129_s;
                stage3_col60[5] = fa_s2_c60_n130_s;
                stage3_col60[6] = fa_s2_c60_n131_s;
                stage3_col60[7] = fa_s2_c60_n132_s;
                stage3_col60[8] = stage2_col60[12];
                stage3_col60[9] = stage2_col60[13];
                stage3_col61[0] = fa_s2_c60_n129_c;
                stage3_col61[1] = fa_s2_c60_n130_c;
                stage3_col61[2] = fa_s2_c60_n131_c;
                stage3_col61[3] = fa_s2_c60_n132_c;
                stage3_col61[4] = fa_s2_c61_n133_s;
                stage3_col61[5] = fa_s2_c61_n134_s;
                stage3_col61[6] = fa_s2_c61_n135_s;
                stage3_col61[7] = fa_s2_c61_n136_s;
                stage3_col61[8] = stage2_col61[12];
                stage3_col61[9] = stage2_col61[13];
                stage3_col62[0] = fa_s2_c61_n133_c;
                stage3_col62[1] = fa_s2_c61_n134_c;
                stage3_col62[2] = fa_s2_c61_n135_c;
                stage3_col62[3] = fa_s2_c61_n136_c;
                stage3_col62[4] = fa_s2_c62_n137_s;
                stage3_col62[5] = fa_s2_c62_n138_s;
                stage3_col62[6] = fa_s2_c62_n139_s;
                stage3_col62[7] = fa_s2_c62_n140_s;
                stage3_col62[8] = stage2_col62[12];
                stage3_col62[9] = stage2_col62[13];
                stage3_col63[0] = fa_s2_c62_n137_c;
                stage3_col63[1] = fa_s2_c62_n138_c;
                stage3_col63[2] = fa_s2_c62_n139_c;
                stage3_col63[3] = fa_s2_c62_n140_c;
                stage3_col63[4] = fa_s2_c63_n141_s;
                stage3_col63[5] = fa_s2_c63_n142_s;
                stage3_col63[6] = fa_s2_c63_n143_s;
                stage3_col63[7] = fa_s2_c63_n144_s;
                stage3_col63[8] = fa_s2_c63_n145_s;
                stage3_col63[9] = stage2_col63[15];
                stage3_col64[0] = fa_s2_c63_n141_c;
                stage3_col64[1] = fa_s2_c63_n142_c;
                stage3_col64[2] = fa_s2_c63_n143_c;
                stage3_col64[3] = fa_s2_c63_n144_c;
                stage3_col64[4] = fa_s2_c63_n145_c;
                stage3_col64[5] = fa_s2_c64_n146_s;
                stage3_col64[6] = fa_s2_c64_n147_s;
                stage3_col64[7] = fa_s2_c64_n148_s;
                stage3_col64[8] = fa_s2_c64_n149_s;
                stage3_col64[9] = stage2_col64[12];
                stage3_col64[10] = stage2_col64[13];
                stage3_col65[0] = fa_s2_c64_n146_c;
                stage3_col65[1] = fa_s2_c64_n147_c;
                stage3_col65[2] = fa_s2_c64_n148_c;
                stage3_col65[3] = fa_s2_c64_n149_c;
                stage3_col65[4] = fa_s2_c65_n150_s;
                stage3_col65[5] = fa_s2_c65_n151_s;
                stage3_col65[6] = fa_s2_c65_n152_s;
                stage3_col65[7] = fa_s2_c65_n153_s;
                stage3_col65[8] = fa_s2_c65_n154_s;
                stage3_col65[9] = stage2_col65[15];
                stage3_col66[0] = fa_s2_c65_n150_c;
                stage3_col66[1] = fa_s2_c65_n151_c;
                stage3_col66[2] = fa_s2_c65_n152_c;
                stage3_col66[3] = fa_s2_c65_n153_c;
                stage3_col66[4] = fa_s2_c65_n154_c;
                stage3_col66[5] = fa_s2_c66_n155_s;
                stage3_col66[6] = fa_s2_c66_n156_s;
                stage3_col66[7] = fa_s2_c66_n157_s;
                stage3_col66[8] = fa_s2_c66_n158_s;
                stage3_col66[9] = stage2_col66[12];
                stage3_col66[10] = stage2_col66[13];
                stage3_col67[0] = fa_s2_c66_n155_c;
                stage3_col67[1] = fa_s2_c66_n156_c;
                stage3_col67[2] = fa_s2_c66_n157_c;
                stage3_col67[3] = fa_s2_c66_n158_c;
                stage3_col67[4] = fa_s2_c67_n159_s;
                stage3_col67[5] = fa_s2_c67_n160_s;
                stage3_col67[6] = fa_s2_c67_n161_s;
                stage3_col67[7] = fa_s2_c67_n162_s;
                stage3_col67[8] = fa_s2_c67_n163_s;
                stage3_col67[9] = stage2_col67[15];
                stage3_col68[0] = fa_s2_c67_n159_c;
                stage3_col68[1] = fa_s2_c67_n160_c;
                stage3_col68[2] = fa_s2_c67_n161_c;
                stage3_col68[3] = fa_s2_c67_n162_c;
                stage3_col68[4] = fa_s2_c67_n163_c;
                stage3_col68[5] = fa_s2_c68_n164_s;
                stage3_col68[6] = fa_s2_c68_n165_s;
                stage3_col68[7] = fa_s2_c68_n166_s;
                stage3_col68[8] = fa_s2_c68_n167_s;
                stage3_col68[9] = stage2_col68[12];
                stage3_col68[10] = stage2_col68[13];
                stage3_col69[0] = fa_s2_c68_n164_c;
                stage3_col69[1] = fa_s2_c68_n165_c;
                stage3_col69[2] = fa_s2_c68_n166_c;
                stage3_col69[3] = fa_s2_c68_n167_c;
                stage3_col69[4] = fa_s2_c69_n168_s;
                stage3_col69[5] = fa_s2_c69_n169_s;
                stage3_col69[6] = fa_s2_c69_n170_s;
                stage3_col69[7] = fa_s2_c69_n171_s;
                stage3_col69[8] = fa_s2_c69_n172_s;
                stage3_col69[9] = stage2_col69[15];
                stage3_col70[0] = fa_s2_c69_n168_c;
                stage3_col70[1] = fa_s2_c69_n169_c;
                stage3_col70[2] = fa_s2_c69_n170_c;
                stage3_col70[3] = fa_s2_c69_n171_c;
                stage3_col70[4] = fa_s2_c69_n172_c;
                stage3_col70[5] = fa_s2_c70_n173_s;
                stage3_col70[6] = fa_s2_c70_n174_s;
                stage3_col70[7] = fa_s2_c70_n175_s;
                stage3_col70[8] = fa_s2_c70_n176_s;
                stage3_col70[9] = stage2_col70[12];
                stage3_col70[10] = stage2_col70[13];
                stage3_col71[0] = fa_s2_c70_n173_c;
                stage3_col71[1] = fa_s2_c70_n174_c;
                stage3_col71[2] = fa_s2_c70_n175_c;
                stage3_col71[3] = fa_s2_c70_n176_c;
                stage3_col71[4] = fa_s2_c71_n177_s;
                stage3_col71[5] = fa_s2_c71_n178_s;
                stage3_col71[6] = fa_s2_c71_n179_s;
                stage3_col71[7] = fa_s2_c71_n180_s;
                stage3_col71[8] = fa_s2_c71_n181_s;
                stage3_col71[9] = stage2_col71[15];
                stage3_col72[0] = fa_s2_c71_n177_c;
                stage3_col72[1] = fa_s2_c71_n178_c;
                stage3_col72[2] = fa_s2_c71_n179_c;
                stage3_col72[3] = fa_s2_c71_n180_c;
                stage3_col72[4] = fa_s2_c71_n181_c;
                stage3_col72[5] = fa_s2_c72_n182_s;
                stage3_col72[6] = fa_s2_c72_n183_s;
                stage3_col72[7] = fa_s2_c72_n184_s;
                stage3_col72[8] = fa_s2_c72_n185_s;
                stage3_col72[9] = stage2_col72[12];
                stage3_col72[10] = stage2_col72[13];
                stage3_col73[0] = fa_s2_c72_n182_c;
                stage3_col73[1] = fa_s2_c72_n183_c;
                stage3_col73[2] = fa_s2_c72_n184_c;
                stage3_col73[3] = fa_s2_c72_n185_c;
                stage3_col73[4] = fa_s2_c73_n186_s;
                stage3_col73[5] = fa_s2_c73_n187_s;
                stage3_col73[6] = fa_s2_c73_n188_s;
                stage3_col73[7] = fa_s2_c73_n189_s;
                stage3_col73[8] = fa_s2_c73_n190_s;
                stage3_col73[9] = stage2_col73[15];
                stage3_col74[0] = fa_s2_c73_n186_c;
                stage3_col74[1] = fa_s2_c73_n187_c;
                stage3_col74[2] = fa_s2_c73_n188_c;
                stage3_col74[3] = fa_s2_c73_n189_c;
                stage3_col74[4] = fa_s2_c73_n190_c;
                stage3_col74[5] = fa_s2_c74_n191_s;
                stage3_col74[6] = fa_s2_c74_n192_s;
                stage3_col74[7] = fa_s2_c74_n193_s;
                stage3_col74[8] = fa_s2_c74_n194_s;
                stage3_col74[9] = stage2_col74[12];
                stage3_col74[10] = stage2_col74[13];
                stage3_col75[0] = fa_s2_c74_n191_c;
                stage3_col75[1] = fa_s2_c74_n192_c;
                stage3_col75[2] = fa_s2_c74_n193_c;
                stage3_col75[3] = fa_s2_c74_n194_c;
                stage3_col75[4] = fa_s2_c75_n195_s;
                stage3_col75[5] = fa_s2_c75_n196_s;
                stage3_col75[6] = fa_s2_c75_n197_s;
                stage3_col75[7] = fa_s2_c75_n198_s;
                stage3_col75[8] = fa_s2_c75_n199_s;
                stage3_col75[9] = stage2_col75[15];
                stage3_col76[0] = fa_s2_c75_n195_c;
                stage3_col76[1] = fa_s2_c75_n196_c;
                stage3_col76[2] = fa_s2_c75_n197_c;
                stage3_col76[3] = fa_s2_c75_n198_c;
                stage3_col76[4] = fa_s2_c75_n199_c;
                stage3_col76[5] = fa_s2_c76_n200_s;
                stage3_col76[6] = fa_s2_c76_n201_s;
                stage3_col76[7] = fa_s2_c76_n202_s;
                stage3_col76[8] = fa_s2_c76_n203_s;
                stage3_col76[9] = stage2_col76[12];
                stage3_col76[10] = stage2_col76[13];
                stage3_col77[0] = fa_s2_c76_n200_c;
                stage3_col77[1] = fa_s2_c76_n201_c;
                stage3_col77[2] = fa_s2_c76_n202_c;
                stage3_col77[3] = fa_s2_c76_n203_c;
                stage3_col77[4] = fa_s2_c77_n204_s;
                stage3_col77[5] = fa_s2_c77_n205_s;
                stage3_col77[6] = fa_s2_c77_n206_s;
                stage3_col77[7] = fa_s2_c77_n207_s;
                stage3_col77[8] = fa_s2_c77_n208_s;
                stage3_col77[9] = stage2_col77[15];
                stage3_col78[0] = fa_s2_c77_n204_c;
                stage3_col78[1] = fa_s2_c77_n205_c;
                stage3_col78[2] = fa_s2_c77_n206_c;
                stage3_col78[3] = fa_s2_c77_n207_c;
                stage3_col78[4] = fa_s2_c77_n208_c;
                stage3_col78[5] = fa_s2_c78_n209_s;
                stage3_col78[6] = fa_s2_c78_n210_s;
                stage3_col78[7] = fa_s2_c78_n211_s;
                stage3_col78[8] = fa_s2_c78_n212_s;
                stage3_col78[9] = stage2_col78[12];
                stage3_col78[10] = stage2_col78[13];
                stage3_col79[0] = fa_s2_c78_n209_c;
                stage3_col79[1] = fa_s2_c78_n210_c;
                stage3_col79[2] = fa_s2_c78_n211_c;
                stage3_col79[3] = fa_s2_c78_n212_c;
                stage3_col79[4] = fa_s2_c79_n213_s;
                stage3_col79[5] = fa_s2_c79_n214_s;
                stage3_col79[6] = fa_s2_c79_n215_s;
                stage3_col79[7] = fa_s2_c79_n216_s;
                stage3_col79[8] = fa_s2_c79_n217_s;
                stage3_col79[9] = stage2_col79[15];
                stage3_col80[0] = fa_s2_c79_n213_c;
                stage3_col80[1] = fa_s2_c79_n214_c;
                stage3_col80[2] = fa_s2_c79_n215_c;
                stage3_col80[3] = fa_s2_c79_n216_c;
                stage3_col80[4] = fa_s2_c79_n217_c;
                stage3_col80[5] = fa_s2_c80_n218_s;
                stage3_col80[6] = fa_s2_c80_n219_s;
                stage3_col80[7] = fa_s2_c80_n220_s;
                stage3_col80[8] = fa_s2_c80_n221_s;
                stage3_col80[9] = stage2_col80[12];
                stage3_col80[10] = stage2_col80[13];
                stage3_col81[0] = fa_s2_c80_n218_c;
                stage3_col81[1] = fa_s2_c80_n219_c;
                stage3_col81[2] = fa_s2_c80_n220_c;
                stage3_col81[3] = fa_s2_c80_n221_c;
                stage3_col81[4] = fa_s2_c81_n222_s;
                stage3_col81[5] = fa_s2_c81_n223_s;
                stage3_col81[6] = fa_s2_c81_n224_s;
                stage3_col81[7] = fa_s2_c81_n225_s;
                stage3_col81[8] = fa_s2_c81_n226_s;
                stage3_col81[9] = stage2_col81[15];
                stage3_col82[0] = fa_s2_c81_n222_c;
                stage3_col82[1] = fa_s2_c81_n223_c;
                stage3_col82[2] = fa_s2_c81_n224_c;
                stage3_col82[3] = fa_s2_c81_n225_c;
                stage3_col82[4] = fa_s2_c81_n226_c;
                stage3_col82[5] = fa_s2_c82_n227_s;
                stage3_col82[6] = fa_s2_c82_n228_s;
                stage3_col82[7] = fa_s2_c82_n229_s;
                stage3_col82[8] = fa_s2_c82_n230_s;
                stage3_col82[9] = stage2_col82[12];
                stage3_col82[10] = stage2_col82[13];
                stage3_col83[0] = fa_s2_c82_n227_c;
                stage3_col83[1] = fa_s2_c82_n228_c;
                stage3_col83[2] = fa_s2_c82_n229_c;
                stage3_col83[3] = fa_s2_c82_n230_c;
                stage3_col83[4] = fa_s2_c83_n231_s;
                stage3_col83[5] = fa_s2_c83_n232_s;
                stage3_col83[6] = fa_s2_c83_n233_s;
                stage3_col83[7] = fa_s2_c83_n234_s;
                stage3_col83[8] = fa_s2_c83_n235_s;
                stage3_col83[9] = stage2_col83[15];
                stage3_col84[0] = fa_s2_c83_n231_c;
                stage3_col84[1] = fa_s2_c83_n232_c;
                stage3_col84[2] = fa_s2_c83_n233_c;
                stage3_col84[3] = fa_s2_c83_n234_c;
                stage3_col84[4] = fa_s2_c83_n235_c;
                stage3_col84[5] = fa_s2_c84_n236_s;
                stage3_col84[6] = fa_s2_c84_n237_s;
                stage3_col84[7] = fa_s2_c84_n238_s;
                stage3_col84[8] = fa_s2_c84_n239_s;
                stage3_col84[9] = stage2_col84[12];
                stage3_col84[10] = stage2_col84[13];
                stage3_col85[0] = fa_s2_c84_n236_c;
                stage3_col85[1] = fa_s2_c84_n237_c;
                stage3_col85[2] = fa_s2_c84_n238_c;
                stage3_col85[3] = fa_s2_c84_n239_c;
                stage3_col85[4] = fa_s2_c85_n240_s;
                stage3_col85[5] = fa_s2_c85_n241_s;
                stage3_col85[6] = fa_s2_c85_n242_s;
                stage3_col85[7] = fa_s2_c85_n243_s;
                stage3_col85[8] = fa_s2_c85_n244_s;
                stage3_col85[9] = stage2_col85[15];
                stage3_col86[0] = fa_s2_c85_n240_c;
                stage3_col86[1] = fa_s2_c85_n241_c;
                stage3_col86[2] = fa_s2_c85_n242_c;
                stage3_col86[3] = fa_s2_c85_n243_c;
                stage3_col86[4] = fa_s2_c85_n244_c;
                stage3_col86[5] = fa_s2_c86_n245_s;
                stage3_col86[6] = fa_s2_c86_n246_s;
                stage3_col86[7] = fa_s2_c86_n247_s;
                stage3_col86[8] = fa_s2_c86_n248_s;
                stage3_col86[9] = stage2_col86[12];
                stage3_col86[10] = stage2_col86[13];
                stage3_col87[0] = fa_s2_c86_n245_c;
                stage3_col87[1] = fa_s2_c86_n246_c;
                stage3_col87[2] = fa_s2_c86_n247_c;
                stage3_col87[3] = fa_s2_c86_n248_c;
                stage3_col87[4] = fa_s2_c87_n249_s;
                stage3_col87[5] = fa_s2_c87_n250_s;
                stage3_col87[6] = fa_s2_c87_n251_s;
                stage3_col87[7] = fa_s2_c87_n252_s;
                stage3_col87[8] = fa_s2_c87_n253_s;
                stage3_col87[9] = stage2_col87[15];
                stage3_col88[0] = fa_s2_c87_n249_c;
                stage3_col88[1] = fa_s2_c87_n250_c;
                stage3_col88[2] = fa_s2_c87_n251_c;
                stage3_col88[3] = fa_s2_c87_n252_c;
                stage3_col88[4] = fa_s2_c87_n253_c;
                stage3_col88[5] = fa_s2_c88_n254_s;
                stage3_col88[6] = fa_s2_c88_n255_s;
                stage3_col88[7] = fa_s2_c88_n256_s;
                stage3_col88[8] = fa_s2_c88_n257_s;
                stage3_col88[9] = stage2_col88[12];
                stage3_col88[10] = stage2_col88[13];
                stage3_col89[0] = fa_s2_c88_n254_c;
                stage3_col89[1] = fa_s2_c88_n255_c;
                stage3_col89[2] = fa_s2_c88_n256_c;
                stage3_col89[3] = fa_s2_c88_n257_c;
                stage3_col89[4] = fa_s2_c89_n258_s;
                stage3_col89[5] = fa_s2_c89_n259_s;
                stage3_col89[6] = fa_s2_c89_n260_s;
                stage3_col89[7] = fa_s2_c89_n261_s;
                stage3_col89[8] = fa_s2_c89_n262_s;
                stage3_col89[9] = stage2_col89[15];
                stage3_col90[0] = fa_s2_c89_n258_c;
                stage3_col90[1] = fa_s2_c89_n259_c;
                stage3_col90[2] = fa_s2_c89_n260_c;
                stage3_col90[3] = fa_s2_c89_n261_c;
                stage3_col90[4] = fa_s2_c89_n262_c;
                stage3_col90[5] = fa_s2_c90_n263_s;
                stage3_col90[6] = fa_s2_c90_n264_s;
                stage3_col90[7] = fa_s2_c90_n265_s;
                stage3_col90[8] = fa_s2_c90_n266_s;
                stage3_col90[9] = stage2_col90[12];
                stage3_col90[10] = stage2_col90[13];
                stage3_col91[0] = fa_s2_c90_n263_c;
                stage3_col91[1] = fa_s2_c90_n264_c;
                stage3_col91[2] = fa_s2_c90_n265_c;
                stage3_col91[3] = fa_s2_c90_n266_c;
                stage3_col91[4] = fa_s2_c91_n267_s;
                stage3_col91[5] = fa_s2_c91_n268_s;
                stage3_col91[6] = fa_s2_c91_n269_s;
                stage3_col91[7] = fa_s2_c91_n270_s;
                stage3_col91[8] = fa_s2_c91_n271_s;
                stage3_col91[9] = stage2_col91[15];
                stage3_col92[0] = fa_s2_c91_n267_c;
                stage3_col92[1] = fa_s2_c91_n268_c;
                stage3_col92[2] = fa_s2_c91_n269_c;
                stage3_col92[3] = fa_s2_c91_n270_c;
                stage3_col92[4] = fa_s2_c91_n271_c;
                stage3_col92[5] = fa_s2_c92_n272_s;
                stage3_col92[6] = fa_s2_c92_n273_s;
                stage3_col92[7] = fa_s2_c92_n274_s;
                stage3_col92[8] = fa_s2_c92_n275_s;
                stage3_col92[9] = stage2_col92[12];
                stage3_col92[10] = stage2_col92[13];
                stage3_col93[0] = fa_s2_c92_n272_c;
                stage3_col93[1] = fa_s2_c92_n273_c;
                stage3_col93[2] = fa_s2_c92_n274_c;
                stage3_col93[3] = fa_s2_c92_n275_c;
                stage3_col93[4] = fa_s2_c93_n276_s;
                stage3_col93[5] = fa_s2_c93_n277_s;
                stage3_col93[6] = fa_s2_c93_n278_s;
                stage3_col93[7] = fa_s2_c93_n279_s;
                stage3_col93[8] = fa_s2_c93_n280_s;
                stage3_col93[9] = stage2_col93[15];
                stage3_col94[0] = fa_s2_c93_n276_c;
                stage3_col94[1] = fa_s2_c93_n277_c;
                stage3_col94[2] = fa_s2_c93_n278_c;
                stage3_col94[3] = fa_s2_c93_n279_c;
                stage3_col94[4] = fa_s2_c93_n280_c;
                stage3_col94[5] = fa_s2_c94_n281_s;
                stage3_col94[6] = fa_s2_c94_n282_s;
                stage3_col94[7] = fa_s2_c94_n283_s;
                stage3_col94[8] = fa_s2_c94_n284_s;
                stage3_col94[9] = stage2_col94[12];
                stage3_col94[10] = stage2_col94[13];
                stage3_col95[0] = fa_s2_c94_n281_c;
                stage3_col95[1] = fa_s2_c94_n282_c;
                stage3_col95[2] = fa_s2_c94_n283_c;
                stage3_col95[3] = fa_s2_c94_n284_c;
                stage3_col95[4] = fa_s2_c95_n285_s;
                stage3_col95[5] = fa_s2_c95_n286_s;
                stage3_col95[6] = fa_s2_c95_n287_s;
                stage3_col95[7] = fa_s2_c95_n288_s;
                stage3_col95[8] = fa_s2_c95_n289_s;
                stage3_col95[9] = stage2_col95[15];
                stage3_col96[0] = fa_s2_c95_n285_c;
                stage3_col96[1] = fa_s2_c95_n286_c;
                stage3_col96[2] = fa_s2_c95_n287_c;
                stage3_col96[3] = fa_s2_c95_n288_c;
                stage3_col96[4] = fa_s2_c95_n289_c;
                stage3_col96[5] = fa_s2_c96_n290_s;
                stage3_col96[6] = fa_s2_c96_n291_s;
                stage3_col96[7] = fa_s2_c96_n292_s;
                stage3_col96[8] = fa_s2_c96_n293_s;
                stage3_col96[9] = stage2_col96[12];
                stage3_col96[10] = stage2_col96[13];
                stage3_col97[0] = fa_s2_c96_n290_c;
                stage3_col97[1] = fa_s2_c96_n291_c;
                stage3_col97[2] = fa_s2_c96_n292_c;
                stage3_col97[3] = fa_s2_c96_n293_c;
                stage3_col97[4] = fa_s2_c97_n294_s;
                stage3_col97[5] = fa_s2_c97_n295_s;
                stage3_col97[6] = fa_s2_c97_n296_s;
                stage3_col97[7] = fa_s2_c97_n297_s;
                stage3_col97[8] = fa_s2_c97_n298_s;
                stage3_col97[9] = stage2_col97[15];
                stage3_col98[0] = fa_s2_c97_n294_c;
                stage3_col98[1] = fa_s2_c97_n295_c;
                stage3_col98[2] = fa_s2_c97_n296_c;
                stage3_col98[3] = fa_s2_c97_n297_c;
                stage3_col98[4] = fa_s2_c97_n298_c;
                stage3_col98[5] = fa_s2_c98_n299_s;
                stage3_col98[6] = fa_s2_c98_n300_s;
                stage3_col98[7] = fa_s2_c98_n301_s;
                stage3_col98[8] = fa_s2_c98_n302_s;
                stage3_col98[9] = stage2_col98[12];
                stage3_col98[10] = stage2_col98[13];
                stage3_col99[0] = fa_s2_c98_n299_c;
                stage3_col99[1] = fa_s2_c98_n300_c;
                stage3_col99[2] = fa_s2_c98_n301_c;
                stage3_col99[3] = fa_s2_c98_n302_c;
                stage3_col99[4] = fa_s2_c99_n303_s;
                stage3_col99[5] = fa_s2_c99_n304_s;
                stage3_col99[6] = fa_s2_c99_n305_s;
                stage3_col99[7] = fa_s2_c99_n306_s;
                stage3_col99[8] = fa_s2_c99_n307_s;
                stage3_col99[9] = stage2_col99[15];
                stage3_col100[0] = fa_s2_c99_n303_c;
                stage3_col100[1] = fa_s2_c99_n304_c;
                stage3_col100[2] = fa_s2_c99_n305_c;
                stage3_col100[3] = fa_s2_c99_n306_c;
                stage3_col100[4] = fa_s2_c99_n307_c;
                stage3_col100[5] = fa_s2_c100_n308_s;
                stage3_col100[6] = fa_s2_c100_n309_s;
                stage3_col100[7] = fa_s2_c100_n310_s;
                stage3_col100[8] = fa_s2_c100_n311_s;
                stage3_col100[9] = stage2_col100[12];
                stage3_col100[10] = stage2_col100[13];
                stage3_col101[0] = fa_s2_c100_n308_c;
                stage3_col101[1] = fa_s2_c100_n309_c;
                stage3_col101[2] = fa_s2_c100_n310_c;
                stage3_col101[3] = fa_s2_c100_n311_c;
                stage3_col101[4] = fa_s2_c101_n312_s;
                stage3_col101[5] = fa_s2_c101_n313_s;
                stage3_col101[6] = fa_s2_c101_n314_s;
                stage3_col101[7] = fa_s2_c101_n315_s;
                stage3_col101[8] = fa_s2_c101_n316_s;
                stage3_col101[9] = stage2_col101[15];
                stage3_col102[0] = fa_s2_c101_n312_c;
                stage3_col102[1] = fa_s2_c101_n313_c;
                stage3_col102[2] = fa_s2_c101_n314_c;
                stage3_col102[3] = fa_s2_c101_n315_c;
                stage3_col102[4] = fa_s2_c101_n316_c;
                stage3_col102[5] = fa_s2_c102_n317_s;
                stage3_col102[6] = fa_s2_c102_n318_s;
                stage3_col102[7] = fa_s2_c102_n319_s;
                stage3_col102[8] = fa_s2_c102_n320_s;
                stage3_col102[9] = stage2_col102[12];
                stage3_col102[10] = stage2_col102[13];
                stage3_col103[0] = fa_s2_c102_n317_c;
                stage3_col103[1] = fa_s2_c102_n318_c;
                stage3_col103[2] = fa_s2_c102_n319_c;
                stage3_col103[3] = fa_s2_c102_n320_c;
                stage3_col103[4] = fa_s2_c103_n321_s;
                stage3_col103[5] = fa_s2_c103_n322_s;
                stage3_col103[6] = fa_s2_c103_n323_s;
                stage3_col103[7] = fa_s2_c103_n324_s;
                stage3_col103[8] = fa_s2_c103_n325_s;
                stage3_col103[9] = stage2_col103[15];
                stage3_col104[0] = fa_s2_c103_n321_c;
                stage3_col104[1] = fa_s2_c103_n322_c;
                stage3_col104[2] = fa_s2_c103_n323_c;
                stage3_col104[3] = fa_s2_c103_n324_c;
                stage3_col104[4] = fa_s2_c103_n325_c;
                stage3_col104[5] = fa_s2_c104_n326_s;
                stage3_col104[6] = fa_s2_c104_n327_s;
                stage3_col104[7] = fa_s2_c104_n328_s;
                stage3_col104[8] = fa_s2_c104_n329_s;
                stage3_col104[9] = stage2_col104[12];
                stage3_col104[10] = stage2_col104[13];
                stage3_col105[0] = fa_s2_c104_n326_c;
                stage3_col105[1] = fa_s2_c104_n327_c;
                stage3_col105[2] = fa_s2_c104_n328_c;
                stage3_col105[3] = fa_s2_c104_n329_c;
                stage3_col105[4] = fa_s2_c105_n330_s;
                stage3_col105[5] = fa_s2_c105_n331_s;
                stage3_col105[6] = fa_s2_c105_n332_s;
                stage3_col105[7] = fa_s2_c105_n333_s;
                stage3_col105[8] = fa_s2_c105_n334_s;
                stage3_col105[9] = stage2_col105[15];
                stage3_col106[0] = fa_s2_c105_n330_c;
                stage3_col106[1] = fa_s2_c105_n331_c;
                stage3_col106[2] = fa_s2_c105_n332_c;
                stage3_col106[3] = fa_s2_c105_n333_c;
                stage3_col106[4] = fa_s2_c105_n334_c;
                stage3_col106[5] = fa_s2_c106_n335_s;
                stage3_col106[6] = fa_s2_c106_n336_s;
                stage3_col106[7] = fa_s2_c106_n337_s;
                stage3_col106[8] = fa_s2_c106_n338_s;
                stage3_col106[9] = stage2_col106[12];
                stage3_col106[10] = stage2_col106[13];
                stage3_col107[0] = fa_s2_c106_n335_c;
                stage3_col107[1] = fa_s2_c106_n336_c;
                stage3_col107[2] = fa_s2_c106_n337_c;
                stage3_col107[3] = fa_s2_c106_n338_c;
                stage3_col107[4] = fa_s2_c107_n339_s;
                stage3_col107[5] = fa_s2_c107_n340_s;
                stage3_col107[6] = fa_s2_c107_n341_s;
                stage3_col107[7] = fa_s2_c107_n342_s;
                stage3_col107[8] = fa_s2_c107_n343_s;
                stage3_col107[9] = stage2_col107[15];
                stage3_col108[0] = fa_s2_c107_n339_c;
                stage3_col108[1] = fa_s2_c107_n340_c;
                stage3_col108[2] = fa_s2_c107_n341_c;
                stage3_col108[3] = fa_s2_c107_n342_c;
                stage3_col108[4] = fa_s2_c107_n343_c;
                stage3_col108[5] = fa_s2_c108_n344_s;
                stage3_col108[6] = fa_s2_c108_n345_s;
                stage3_col108[7] = fa_s2_c108_n346_s;
                stage3_col108[8] = fa_s2_c108_n347_s;
                stage3_col108[9] = stage2_col108[12];
                stage3_col108[10] = stage2_col108[13];
                stage3_col109[0] = fa_s2_c108_n344_c;
                stage3_col109[1] = fa_s2_c108_n345_c;
                stage3_col109[2] = fa_s2_c108_n346_c;
                stage3_col109[3] = fa_s2_c108_n347_c;
                stage3_col109[4] = fa_s2_c109_n348_s;
                stage3_col109[5] = fa_s2_c109_n349_s;
                stage3_col109[6] = fa_s2_c109_n350_s;
                stage3_col109[7] = fa_s2_c109_n351_s;
                stage3_col109[8] = fa_s2_c109_n352_s;
                stage3_col109[9] = stage2_col109[15];
                stage3_col110[0] = fa_s2_c109_n348_c;
                stage3_col110[1] = fa_s2_c109_n349_c;
                stage3_col110[2] = fa_s2_c109_n350_c;
                stage3_col110[3] = fa_s2_c109_n351_c;
                stage3_col110[4] = fa_s2_c109_n352_c;
                stage3_col110[5] = fa_s2_c110_n353_s;
                stage3_col110[6] = fa_s2_c110_n354_s;
                stage3_col110[7] = fa_s2_c110_n355_s;
                stage3_col110[8] = fa_s2_c110_n356_s;
                stage3_col110[9] = stage2_col110[12];
                stage3_col110[10] = stage2_col110[13];
                stage3_col111[0] = fa_s2_c110_n353_c;
                stage3_col111[1] = fa_s2_c110_n354_c;
                stage3_col111[2] = fa_s2_c110_n355_c;
                stage3_col111[3] = fa_s2_c110_n356_c;
                stage3_col111[4] = fa_s2_c111_n357_s;
                stage3_col111[5] = fa_s2_c111_n358_s;
                stage3_col111[6] = fa_s2_c111_n359_s;
                stage3_col111[7] = fa_s2_c111_n360_s;
                stage3_col111[8] = fa_s2_c111_n361_s;
                stage3_col111[9] = stage2_col111[15];
                stage3_col112[0] = fa_s2_c111_n357_c;
                stage3_col112[1] = fa_s2_c111_n358_c;
                stage3_col112[2] = fa_s2_c111_n359_c;
                stage3_col112[3] = fa_s2_c111_n360_c;
                stage3_col112[4] = fa_s2_c111_n361_c;
                stage3_col112[5] = fa_s2_c112_n362_s;
                stage3_col112[6] = fa_s2_c112_n363_s;
                stage3_col112[7] = fa_s2_c112_n364_s;
                stage3_col112[8] = fa_s2_c112_n365_s;
                stage3_col112[9] = stage2_col112[12];
                stage3_col112[10] = stage2_col112[13];
                stage3_col113[0] = fa_s2_c112_n362_c;
                stage3_col113[1] = fa_s2_c112_n363_c;
                stage3_col113[2] = fa_s2_c112_n364_c;
                stage3_col113[3] = fa_s2_c112_n365_c;
                stage3_col113[4] = fa_s2_c113_n366_s;
                stage3_col113[5] = fa_s2_c113_n367_s;
                stage3_col113[6] = fa_s2_c113_n368_s;
                stage3_col113[7] = fa_s2_c113_n369_s;
                stage3_col113[8] = fa_s2_c113_n370_s;
                stage3_col113[9] = stage2_col113[15];
                stage3_col114[0] = fa_s2_c113_n366_c;
                stage3_col114[1] = fa_s2_c113_n367_c;
                stage3_col114[2] = fa_s2_c113_n368_c;
                stage3_col114[3] = fa_s2_c113_n369_c;
                stage3_col114[4] = fa_s2_c113_n370_c;
                stage3_col114[5] = fa_s2_c114_n371_s;
                stage3_col114[6] = fa_s2_c114_n372_s;
                stage3_col114[7] = fa_s2_c114_n373_s;
                stage3_col114[8] = fa_s2_c114_n374_s;
                stage3_col114[9] = stage2_col114[12];
                stage3_col114[10] = stage2_col114[13];
                stage3_col115[0] = fa_s2_c114_n371_c;
                stage3_col115[1] = fa_s2_c114_n372_c;
                stage3_col115[2] = fa_s2_c114_n373_c;
                stage3_col115[3] = fa_s2_c114_n374_c;
                stage3_col115[4] = fa_s2_c115_n375_s;
                stage3_col115[5] = fa_s2_c115_n376_s;
                stage3_col115[6] = fa_s2_c115_n377_s;
                stage3_col115[7] = fa_s2_c115_n378_s;
                stage3_col115[8] = fa_s2_c115_n379_s;
                stage3_col115[9] = stage2_col115[15];
                stage3_col116[0] = fa_s2_c115_n375_c;
                stage3_col116[1] = fa_s2_c115_n376_c;
                stage3_col116[2] = fa_s2_c115_n377_c;
                stage3_col116[3] = fa_s2_c115_n378_c;
                stage3_col116[4] = fa_s2_c115_n379_c;
                stage3_col116[5] = fa_s2_c116_n380_s;
                stage3_col116[6] = fa_s2_c116_n381_s;
                stage3_col116[7] = fa_s2_c116_n382_s;
                stage3_col116[8] = fa_s2_c116_n383_s;
                stage3_col116[9] = stage2_col116[12];
                stage3_col116[10] = stage2_col116[13];
                stage3_col117[0] = fa_s2_c116_n380_c;
                stage3_col117[1] = fa_s2_c116_n381_c;
                stage3_col117[2] = fa_s2_c116_n382_c;
                stage3_col117[3] = fa_s2_c116_n383_c;
                stage3_col117[4] = fa_s2_c117_n384_s;
                stage3_col117[5] = fa_s2_c117_n385_s;
                stage3_col117[6] = fa_s2_c117_n386_s;
                stage3_col117[7] = fa_s2_c117_n387_s;
                stage3_col117[8] = fa_s2_c117_n388_s;
                stage3_col117[9] = stage2_col117[15];
                stage3_col118[0] = fa_s2_c117_n384_c;
                stage3_col118[1] = fa_s2_c117_n385_c;
                stage3_col118[2] = fa_s2_c117_n386_c;
                stage3_col118[3] = fa_s2_c117_n387_c;
                stage3_col118[4] = fa_s2_c117_n388_c;
                stage3_col118[5] = fa_s2_c118_n389_s;
                stage3_col118[6] = fa_s2_c118_n390_s;
                stage3_col118[7] = fa_s2_c118_n391_s;
                stage3_col118[8] = fa_s2_c118_n392_s;
                stage3_col118[9] = stage2_col118[12];
                stage3_col118[10] = stage2_col118[13];
                stage3_col119[0] = fa_s2_c118_n389_c;
                stage3_col119[1] = fa_s2_c118_n390_c;
                stage3_col119[2] = fa_s2_c118_n391_c;
                stage3_col119[3] = fa_s2_c118_n392_c;
                stage3_col119[4] = fa_s2_c119_n393_s;
                stage3_col119[5] = fa_s2_c119_n394_s;
                stage3_col119[6] = fa_s2_c119_n395_s;
                stage3_col119[7] = fa_s2_c119_n396_s;
                stage3_col119[8] = fa_s2_c119_n397_s;
                stage3_col119[9] = stage2_col119[15];
                stage3_col120[0] = fa_s2_c119_n393_c;
                stage3_col120[1] = fa_s2_c119_n394_c;
                stage3_col120[2] = fa_s2_c119_n395_c;
                stage3_col120[3] = fa_s2_c119_n396_c;
                stage3_col120[4] = fa_s2_c119_n397_c;
                stage3_col120[5] = fa_s2_c120_n398_s;
                stage3_col120[6] = fa_s2_c120_n399_s;
                stage3_col120[7] = fa_s2_c120_n400_s;
                stage3_col120[8] = fa_s2_c120_n401_s;
                stage3_col120[9] = stage2_col120[12];
                stage3_col120[10] = stage2_col120[13];
                stage3_col121[0] = fa_s2_c120_n398_c;
                stage3_col121[1] = fa_s2_c120_n399_c;
                stage3_col121[2] = fa_s2_c120_n400_c;
                stage3_col121[3] = fa_s2_c120_n401_c;
                stage3_col121[4] = fa_s2_c121_n402_s;
                stage3_col121[5] = fa_s2_c121_n403_s;
                stage3_col121[6] = fa_s2_c121_n404_s;
                stage3_col121[7] = fa_s2_c121_n405_s;
                stage3_col121[8] = fa_s2_c121_n406_s;
                stage3_col121[9] = stage2_col121[15];
                stage3_col122[0] = fa_s2_c121_n402_c;
                stage3_col122[1] = fa_s2_c121_n403_c;
                stage3_col122[2] = fa_s2_c121_n404_c;
                stage3_col122[3] = fa_s2_c121_n405_c;
                stage3_col122[4] = fa_s2_c121_n406_c;
                stage3_col122[5] = fa_s2_c122_n407_s;
                stage3_col122[6] = fa_s2_c122_n408_s;
                stage3_col122[7] = fa_s2_c122_n409_s;
                stage3_col122[8] = fa_s2_c122_n410_s;
                stage3_col122[9] = stage2_col122[12];
                stage3_col122[10] = stage2_col122[13];
                stage3_col123[0] = fa_s2_c122_n407_c;
                stage3_col123[1] = fa_s2_c122_n408_c;
                stage3_col123[2] = fa_s2_c122_n409_c;
                stage3_col123[3] = fa_s2_c122_n410_c;
                stage3_col123[4] = fa_s2_c123_n411_s;
                stage3_col123[5] = fa_s2_c123_n412_s;
                stage3_col123[6] = fa_s2_c123_n413_s;
                stage3_col123[7] = fa_s2_c123_n414_s;
                stage3_col123[8] = fa_s2_c123_n415_s;
                stage3_col123[9] = stage2_col123[15];
                stage3_col124[0] = fa_s2_c123_n411_c;
                stage3_col124[1] = fa_s2_c123_n412_c;
                stage3_col124[2] = fa_s2_c123_n413_c;
                stage3_col124[3] = fa_s2_c123_n414_c;
                stage3_col124[4] = fa_s2_c123_n415_c;
                stage3_col124[5] = fa_s2_c124_n416_s;
                stage3_col124[6] = fa_s2_c124_n417_s;
                stage3_col124[7] = fa_s2_c124_n418_s;
                stage3_col124[8] = fa_s2_c124_n419_s;
                stage3_col124[9] = stage2_col124[12];
                stage3_col124[10] = stage2_col124[13];
                stage3_col125[0] = fa_s2_c124_n416_c;
                stage3_col125[1] = fa_s2_c124_n417_c;
                stage3_col125[2] = fa_s2_c124_n418_c;
                stage3_col125[3] = fa_s2_c124_n419_c;
                stage3_col125[4] = fa_s2_c125_n420_s;
                stage3_col125[5] = fa_s2_c125_n421_s;
                stage3_col125[6] = fa_s2_c125_n422_s;
                stage3_col125[7] = fa_s2_c125_n423_s;
                stage3_col125[8] = fa_s2_c125_n424_s;
                stage3_col125[9] = stage2_col125[15];
                stage3_col126[0] = fa_s2_c125_n420_c;
                stage3_col126[1] = fa_s2_c125_n421_c;
                stage3_col126[2] = fa_s2_c125_n422_c;
                stage3_col126[3] = fa_s2_c125_n423_c;
                stage3_col126[4] = fa_s2_c125_n424_c;
                stage3_col126[5] = fa_s2_c126_n425_s;
                stage3_col126[6] = fa_s2_c126_n426_s;
                stage3_col126[7] = fa_s2_c126_n427_s;
                stage3_col126[8] = fa_s2_c126_n428_s;
                stage3_col126[9] = stage2_col126[12];
                stage3_col126[10] = stage2_col126[13];
                stage3_col127[0] = fa_s2_c126_n425_c;
                stage3_col127[1] = fa_s2_c126_n426_c;
                stage3_col127[2] = fa_s2_c126_n427_c;
                stage3_col127[3] = fa_s2_c126_n428_c;
                stage3_col127[4] = stage2_col127[0];
                stage3_col127[5] = stage2_col127[1];
                stage3_col127[6] = stage2_col127[2];
                stage3_col127[7] = stage2_col127[3];
                stage3_col127[8] = stage2_col127[4];
                stage3_col127[9] = stage2_col127[5];
                stage3_col127[10] = stage2_col127[6];
                stage3_col127[11] = stage2_col127[7];
                stage3_col127[12] = stage2_col127[8];
                stage3_col127[13] = stage2_col127[9];
                stage3_col127[14] = stage2_col127[10];
                stage3_col127[15] = stage2_col127[11];
                stage3_col127[16] = stage2_col127[12];
                stage3_col127[17] = stage2_col127[13];
                stage3_col127[18] = stage2_col127[14];
                stage3_col127[19] = stage2_col127[15];
                stage3_col127[20] = stage2_col127[16];
                stage3_col127[21] = stage2_col127[17];
                stage3_col127[22] = stage2_col127[18];
                stage3_col127[23] = stage2_col127[18];
                stage3_col127[24] = stage2_col127[18];
                stage3_col127[25] = stage2_col127[18];
                stage3_col127[26] = stage2_col127[18];
                stage3_col127[27] = stage2_col127[18];
                stage3_col127[28] = stage2_col127[18];
                stage3_col127[29] = stage2_col127[18];
                stage3_col127[30] = stage2_col127[18];
                stage3_col127[31] = stage2_col127[18];
                stage3_col127[32] = stage2_col127[18];
                stage3_col127[33] = stage2_col127[18];
                stage3_col127[34] = stage2_col127[18];
                stage3_col127[35] = stage2_col127[18];
                stage3_col127[36] = stage2_col127[18];
                stage3_col127[37] = stage2_col127[18];
                stage3_col127[38] = stage2_col127[18];
                stage3_col127[39] = stage2_col127[18];
                stage3_col127[40] = stage2_col127[18];
                stage3_col127[41] = stage2_col127[18];
                stage3_col127[42] = stage2_col127[18];
                stage3_col127[43] = stage2_col127[18];
                stage3_col127[44] = stage2_col127[18];
                stage3_col127[45] = stage2_col127[18];
                stage3_col127[46] = stage2_col127[18];
                stage3_col127[47] = stage2_col127[18];
                stage3_col127[48] = stage2_col127[18];
                stage3_col127[49] = stage2_col127[18];
                stage3_col127[50] = stage2_col127[18];
                stage3_col127[51] = stage2_col127[18];
                stage3_col127[52] = stage2_col127[18];
                stage3_col127[53] = stage2_col127[18];
            end
        end
    endgenerate

    // Stage 4: Reduction
    fa fa_s3_c5_n0 (
        .a(stage3_col5[0]),
        .b(stage3_col5[1]),
        .c_in(stage3_col5[2]),
        .s(fa_s3_c5_n0_s),
        .c_out(fa_s3_c5_n0_c)
    );

    fa fa_s3_c13_n1 (
        .a(stage3_col13[0]),
        .b(stage3_col13[1]),
        .c_in(stage3_col13[2]),
        .s(fa_s3_c13_n1_s),
        .c_out(fa_s3_c13_n1_c)
    );

    fa fa_s3_c14_n2 (
        .a(stage3_col14[0]),
        .b(stage3_col14[1]),
        .c_in(stage3_col14[2]),
        .s(fa_s3_c14_n2_s),
        .c_out(fa_s3_c14_n2_c)
    );

    fa fa_s3_c15_n3 (
        .a(stage3_col15[0]),
        .b(stage3_col15[1]),
        .c_in(stage3_col15[2]),
        .s(fa_s3_c15_n3_s),
        .c_out(fa_s3_c15_n3_c)
    );

    fa fa_s3_c16_n4 (
        .a(stage3_col16[0]),
        .b(stage3_col16[1]),
        .c_in(stage3_col16[2]),
        .s(fa_s3_c16_n4_s),
        .c_out(fa_s3_c16_n4_c)
    );

    fa fa_s3_c17_n5 (
        .a(stage3_col17[0]),
        .b(stage3_col17[1]),
        .c_in(stage3_col17[2]),
        .s(fa_s3_c17_n5_s),
        .c_out(fa_s3_c17_n5_c)
    );

    fa fa_s3_c18_n6 (
        .a(stage3_col18[0]),
        .b(stage3_col18[1]),
        .c_in(stage3_col18[2]),
        .s(fa_s3_c18_n6_s),
        .c_out(fa_s3_c18_n6_c)
    );

    fa fa_s3_c19_n7 (
        .a(stage3_col19[0]),
        .b(stage3_col19[1]),
        .c_in(stage3_col19[2]),
        .s(fa_s3_c19_n7_s),
        .c_out(fa_s3_c19_n7_c)
    );

    fa fa_s3_c20_n8 (
        .a(stage3_col20[0]),
        .b(stage3_col20[1]),
        .c_in(stage3_col20[2]),
        .s(fa_s3_c20_n8_s),
        .c_out(fa_s3_c20_n8_c)
    );

    fa fa_s3_c21_n9 (
        .a(stage3_col21[0]),
        .b(stage3_col21[1]),
        .c_in(stage3_col21[2]),
        .s(fa_s3_c21_n9_s),
        .c_out(fa_s3_c21_n9_c)
    );

    fa fa_s3_c22_n10 (
        .a(stage3_col22[0]),
        .b(stage3_col22[1]),
        .c_in(stage3_col22[2]),
        .s(fa_s3_c22_n10_s),
        .c_out(fa_s3_c22_n10_c)
    );

    fa fa_s3_c23_n11 (
        .a(stage3_col23[0]),
        .b(stage3_col23[1]),
        .c_in(stage3_col23[2]),
        .s(fa_s3_c23_n11_s),
        .c_out(fa_s3_c23_n11_c)
    );

    fa fa_s3_c24_n12 (
        .a(stage3_col24[0]),
        .b(stage3_col24[1]),
        .c_in(stage3_col24[2]),
        .s(fa_s3_c24_n12_s),
        .c_out(fa_s3_c24_n12_c)
    );

    fa fa_s3_c25_n13 (
        .a(stage3_col25[0]),
        .b(stage3_col25[1]),
        .c_in(stage3_col25[2]),
        .s(fa_s3_c25_n13_s),
        .c_out(fa_s3_c25_n13_c)
    );

    fa fa_s3_c26_n14 (
        .a(stage3_col26[0]),
        .b(stage3_col26[1]),
        .c_in(stage3_col26[2]),
        .s(fa_s3_c26_n14_s),
        .c_out(fa_s3_c26_n14_c)
    );

    fa fa_s3_c27_n15 (
        .a(stage3_col27[0]),
        .b(stage3_col27[1]),
        .c_in(stage3_col27[2]),
        .s(fa_s3_c27_n15_s),
        .c_out(fa_s3_c27_n15_c)
    );

    fa fa_s3_c27_n16 (
        .a(stage3_col27[3]),
        .b(stage3_col27[4]),
        .c_in(stage3_col27[5]),
        .s(fa_s3_c27_n16_s),
        .c_out(fa_s3_c27_n16_c)
    );

    fa fa_s3_c28_n17 (
        .a(stage3_col28[0]),
        .b(stage3_col28[1]),
        .c_in(stage3_col28[2]),
        .s(fa_s3_c28_n17_s),
        .c_out(fa_s3_c28_n17_c)
    );

    fa fa_s3_c29_n18 (
        .a(stage3_col29[0]),
        .b(stage3_col29[1]),
        .c_in(stage3_col29[2]),
        .s(fa_s3_c29_n18_s),
        .c_out(fa_s3_c29_n18_c)
    );

    fa fa_s3_c30_n19 (
        .a(stage3_col30[0]),
        .b(stage3_col30[1]),
        .c_in(stage3_col30[2]),
        .s(fa_s3_c30_n19_s),
        .c_out(fa_s3_c30_n19_c)
    );

    fa fa_s3_c31_n20 (
        .a(stage3_col31[0]),
        .b(stage3_col31[1]),
        .c_in(stage3_col31[2]),
        .s(fa_s3_c31_n20_s),
        .c_out(fa_s3_c31_n20_c)
    );

    fa fa_s3_c32_n21 (
        .a(stage3_col32[0]),
        .b(stage3_col32[1]),
        .c_in(stage3_col32[2]),
        .s(fa_s3_c32_n21_s),
        .c_out(fa_s3_c32_n21_c)
    );

    fa fa_s3_c32_n22 (
        .a(stage3_col32[3]),
        .b(stage3_col32[4]),
        .c_in(stage3_col32[5]),
        .s(fa_s3_c32_n22_s),
        .c_out(fa_s3_c32_n22_c)
    );

    fa fa_s3_c33_n23 (
        .a(stage3_col33[0]),
        .b(stage3_col33[1]),
        .c_in(stage3_col33[2]),
        .s(fa_s3_c33_n23_s),
        .c_out(fa_s3_c33_n23_c)
    );

    fa fa_s3_c33_n24 (
        .a(stage3_col33[3]),
        .b(stage3_col33[4]),
        .c_in(stage3_col33[5]),
        .s(fa_s3_c33_n24_s),
        .c_out(fa_s3_c33_n24_c)
    );

    fa fa_s3_c34_n25 (
        .a(stage3_col34[0]),
        .b(stage3_col34[1]),
        .c_in(stage3_col34[2]),
        .s(fa_s3_c34_n25_s),
        .c_out(fa_s3_c34_n25_c)
    );

    fa fa_s3_c34_n26 (
        .a(stage3_col34[3]),
        .b(stage3_col34[4]),
        .c_in(stage3_col34[5]),
        .s(fa_s3_c34_n26_s),
        .c_out(fa_s3_c34_n26_c)
    );

    fa fa_s3_c35_n27 (
        .a(stage3_col35[0]),
        .b(stage3_col35[1]),
        .c_in(stage3_col35[2]),
        .s(fa_s3_c35_n27_s),
        .c_out(fa_s3_c35_n27_c)
    );

    fa fa_s3_c35_n28 (
        .a(stage3_col35[3]),
        .b(stage3_col35[4]),
        .c_in(stage3_col35[5]),
        .s(fa_s3_c35_n28_s),
        .c_out(fa_s3_c35_n28_c)
    );

    fa fa_s3_c36_n29 (
        .a(stage3_col36[0]),
        .b(stage3_col36[1]),
        .c_in(stage3_col36[2]),
        .s(fa_s3_c36_n29_s),
        .c_out(fa_s3_c36_n29_c)
    );

    fa fa_s3_c36_n30 (
        .a(stage3_col36[3]),
        .b(stage3_col36[4]),
        .c_in(stage3_col36[5]),
        .s(fa_s3_c36_n30_s),
        .c_out(fa_s3_c36_n30_c)
    );

    fa fa_s3_c37_n31 (
        .a(stage3_col37[0]),
        .b(stage3_col37[1]),
        .c_in(stage3_col37[2]),
        .s(fa_s3_c37_n31_s),
        .c_out(fa_s3_c37_n31_c)
    );

    fa fa_s3_c37_n32 (
        .a(stage3_col37[3]),
        .b(stage3_col37[4]),
        .c_in(stage3_col37[5]),
        .s(fa_s3_c37_n32_s),
        .c_out(fa_s3_c37_n32_c)
    );

    fa fa_s3_c38_n33 (
        .a(stage3_col38[0]),
        .b(stage3_col38[1]),
        .c_in(stage3_col38[2]),
        .s(fa_s3_c38_n33_s),
        .c_out(fa_s3_c38_n33_c)
    );

    fa fa_s3_c38_n34 (
        .a(stage3_col38[3]),
        .b(stage3_col38[4]),
        .c_in(stage3_col38[5]),
        .s(fa_s3_c38_n34_s),
        .c_out(fa_s3_c38_n34_c)
    );

    fa fa_s3_c39_n35 (
        .a(stage3_col39[0]),
        .b(stage3_col39[1]),
        .c_in(stage3_col39[2]),
        .s(fa_s3_c39_n35_s),
        .c_out(fa_s3_c39_n35_c)
    );

    fa fa_s3_c39_n36 (
        .a(stage3_col39[3]),
        .b(stage3_col39[4]),
        .c_in(stage3_col39[5]),
        .s(fa_s3_c39_n36_s),
        .c_out(fa_s3_c39_n36_c)
    );

    fa fa_s3_c40_n37 (
        .a(stage3_col40[0]),
        .b(stage3_col40[1]),
        .c_in(stage3_col40[2]),
        .s(fa_s3_c40_n37_s),
        .c_out(fa_s3_c40_n37_c)
    );

    fa fa_s3_c40_n38 (
        .a(stage3_col40[3]),
        .b(stage3_col40[4]),
        .c_in(stage3_col40[5]),
        .s(fa_s3_c40_n38_s),
        .c_out(fa_s3_c40_n38_c)
    );

    fa fa_s3_c41_n39 (
        .a(stage3_col41[0]),
        .b(stage3_col41[1]),
        .c_in(stage3_col41[2]),
        .s(fa_s3_c41_n39_s),
        .c_out(fa_s3_c41_n39_c)
    );

    fa fa_s3_c41_n40 (
        .a(stage3_col41[3]),
        .b(stage3_col41[4]),
        .c_in(stage3_col41[5]),
        .s(fa_s3_c41_n40_s),
        .c_out(fa_s3_c41_n40_c)
    );

    fa fa_s3_c42_n41 (
        .a(stage3_col42[0]),
        .b(stage3_col42[1]),
        .c_in(stage3_col42[2]),
        .s(fa_s3_c42_n41_s),
        .c_out(fa_s3_c42_n41_c)
    );

    fa fa_s3_c42_n42 (
        .a(stage3_col42[3]),
        .b(stage3_col42[4]),
        .c_in(stage3_col42[5]),
        .s(fa_s3_c42_n42_s),
        .c_out(fa_s3_c42_n42_c)
    );

    fa fa_s3_c43_n43 (
        .a(stage3_col43[0]),
        .b(stage3_col43[1]),
        .c_in(stage3_col43[2]),
        .s(fa_s3_c43_n43_s),
        .c_out(fa_s3_c43_n43_c)
    );

    fa fa_s3_c43_n44 (
        .a(stage3_col43[3]),
        .b(stage3_col43[4]),
        .c_in(stage3_col43[5]),
        .s(fa_s3_c43_n44_s),
        .c_out(fa_s3_c43_n44_c)
    );

    fa fa_s3_c44_n45 (
        .a(stage3_col44[0]),
        .b(stage3_col44[1]),
        .c_in(stage3_col44[2]),
        .s(fa_s3_c44_n45_s),
        .c_out(fa_s3_c44_n45_c)
    );

    fa fa_s3_c44_n46 (
        .a(stage3_col44[3]),
        .b(stage3_col44[4]),
        .c_in(stage3_col44[5]),
        .s(fa_s3_c44_n46_s),
        .c_out(fa_s3_c44_n46_c)
    );

    fa fa_s3_c45_n47 (
        .a(stage3_col45[0]),
        .b(stage3_col45[1]),
        .c_in(stage3_col45[2]),
        .s(fa_s3_c45_n47_s),
        .c_out(fa_s3_c45_n47_c)
    );

    fa fa_s3_c45_n48 (
        .a(stage3_col45[3]),
        .b(stage3_col45[4]),
        .c_in(stage3_col45[5]),
        .s(fa_s3_c45_n48_s),
        .c_out(fa_s3_c45_n48_c)
    );

    fa fa_s3_c46_n49 (
        .a(stage3_col46[0]),
        .b(stage3_col46[1]),
        .c_in(stage3_col46[2]),
        .s(fa_s3_c46_n49_s),
        .c_out(fa_s3_c46_n49_c)
    );

    fa fa_s3_c46_n50 (
        .a(stage3_col46[3]),
        .b(stage3_col46[4]),
        .c_in(stage3_col46[5]),
        .s(fa_s3_c46_n50_s),
        .c_out(fa_s3_c46_n50_c)
    );

    fa fa_s3_c46_n51 (
        .a(stage3_col46[6]),
        .b(stage3_col46[7]),
        .c_in(stage3_col46[8]),
        .s(fa_s3_c46_n51_s),
        .c_out(fa_s3_c46_n51_c)
    );

    fa fa_s3_c47_n52 (
        .a(stage3_col47[0]),
        .b(stage3_col47[1]),
        .c_in(stage3_col47[2]),
        .s(fa_s3_c47_n52_s),
        .c_out(fa_s3_c47_n52_c)
    );

    fa fa_s3_c47_n53 (
        .a(stage3_col47[3]),
        .b(stage3_col47[4]),
        .c_in(stage3_col47[5]),
        .s(fa_s3_c47_n53_s),
        .c_out(fa_s3_c47_n53_c)
    );

    fa fa_s3_c48_n54 (
        .a(stage3_col48[0]),
        .b(stage3_col48[1]),
        .c_in(stage3_col48[2]),
        .s(fa_s3_c48_n54_s),
        .c_out(fa_s3_c48_n54_c)
    );

    fa fa_s3_c48_n55 (
        .a(stage3_col48[3]),
        .b(stage3_col48[4]),
        .c_in(stage3_col48[5]),
        .s(fa_s3_c48_n55_s),
        .c_out(fa_s3_c48_n55_c)
    );

    fa fa_s3_c49_n56 (
        .a(stage3_col49[0]),
        .b(stage3_col49[1]),
        .c_in(stage3_col49[2]),
        .s(fa_s3_c49_n56_s),
        .c_out(fa_s3_c49_n56_c)
    );

    fa fa_s3_c49_n57 (
        .a(stage3_col49[3]),
        .b(stage3_col49[4]),
        .c_in(stage3_col49[5]),
        .s(fa_s3_c49_n57_s),
        .c_out(fa_s3_c49_n57_c)
    );

    fa fa_s3_c50_n58 (
        .a(stage3_col50[0]),
        .b(stage3_col50[1]),
        .c_in(stage3_col50[2]),
        .s(fa_s3_c50_n58_s),
        .c_out(fa_s3_c50_n58_c)
    );

    fa fa_s3_c50_n59 (
        .a(stage3_col50[3]),
        .b(stage3_col50[4]),
        .c_in(stage3_col50[5]),
        .s(fa_s3_c50_n59_s),
        .c_out(fa_s3_c50_n59_c)
    );

    fa fa_s3_c51_n60 (
        .a(stage3_col51[0]),
        .b(stage3_col51[1]),
        .c_in(stage3_col51[2]),
        .s(fa_s3_c51_n60_s),
        .c_out(fa_s3_c51_n60_c)
    );

    fa fa_s3_c51_n61 (
        .a(stage3_col51[3]),
        .b(stage3_col51[4]),
        .c_in(stage3_col51[5]),
        .s(fa_s3_c51_n61_s),
        .c_out(fa_s3_c51_n61_c)
    );

    fa fa_s3_c52_n62 (
        .a(stage3_col52[0]),
        .b(stage3_col52[1]),
        .c_in(stage3_col52[2]),
        .s(fa_s3_c52_n62_s),
        .c_out(fa_s3_c52_n62_c)
    );

    fa fa_s3_c52_n63 (
        .a(stage3_col52[3]),
        .b(stage3_col52[4]),
        .c_in(stage3_col52[5]),
        .s(fa_s3_c52_n63_s),
        .c_out(fa_s3_c52_n63_c)
    );

    fa fa_s3_c53_n64 (
        .a(stage3_col53[0]),
        .b(stage3_col53[1]),
        .c_in(stage3_col53[2]),
        .s(fa_s3_c53_n64_s),
        .c_out(fa_s3_c53_n64_c)
    );

    fa fa_s3_c53_n65 (
        .a(stage3_col53[3]),
        .b(stage3_col53[4]),
        .c_in(stage3_col53[5]),
        .s(fa_s3_c53_n65_s),
        .c_out(fa_s3_c53_n65_c)
    );

    fa fa_s3_c54_n66 (
        .a(stage3_col54[0]),
        .b(stage3_col54[1]),
        .c_in(stage3_col54[2]),
        .s(fa_s3_c54_n66_s),
        .c_out(fa_s3_c54_n66_c)
    );

    fa fa_s3_c54_n67 (
        .a(stage3_col54[3]),
        .b(stage3_col54[4]),
        .c_in(stage3_col54[5]),
        .s(fa_s3_c54_n67_s),
        .c_out(fa_s3_c54_n67_c)
    );

    fa fa_s3_c54_n68 (
        .a(stage3_col54[6]),
        .b(stage3_col54[7]),
        .c_in(stage3_col54[8]),
        .s(fa_s3_c54_n68_s),
        .c_out(fa_s3_c54_n68_c)
    );

    fa fa_s3_c55_n69 (
        .a(stage3_col55[0]),
        .b(stage3_col55[1]),
        .c_in(stage3_col55[2]),
        .s(fa_s3_c55_n69_s),
        .c_out(fa_s3_c55_n69_c)
    );

    fa fa_s3_c55_n70 (
        .a(stage3_col55[3]),
        .b(stage3_col55[4]),
        .c_in(stage3_col55[5]),
        .s(fa_s3_c55_n70_s),
        .c_out(fa_s3_c55_n70_c)
    );

    fa fa_s3_c55_n71 (
        .a(stage3_col55[6]),
        .b(stage3_col55[7]),
        .c_in(stage3_col55[8]),
        .s(fa_s3_c55_n71_s),
        .c_out(fa_s3_c55_n71_c)
    );

    fa fa_s3_c56_n72 (
        .a(stage3_col56[0]),
        .b(stage3_col56[1]),
        .c_in(stage3_col56[2]),
        .s(fa_s3_c56_n72_s),
        .c_out(fa_s3_c56_n72_c)
    );

    fa fa_s3_c56_n73 (
        .a(stage3_col56[3]),
        .b(stage3_col56[4]),
        .c_in(stage3_col56[5]),
        .s(fa_s3_c56_n73_s),
        .c_out(fa_s3_c56_n73_c)
    );

    fa fa_s3_c56_n74 (
        .a(stage3_col56[6]),
        .b(stage3_col56[7]),
        .c_in(stage3_col56[8]),
        .s(fa_s3_c56_n74_s),
        .c_out(fa_s3_c56_n74_c)
    );

    fa fa_s3_c57_n75 (
        .a(stage3_col57[0]),
        .b(stage3_col57[1]),
        .c_in(stage3_col57[2]),
        .s(fa_s3_c57_n75_s),
        .c_out(fa_s3_c57_n75_c)
    );

    fa fa_s3_c57_n76 (
        .a(stage3_col57[3]),
        .b(stage3_col57[4]),
        .c_in(stage3_col57[5]),
        .s(fa_s3_c57_n76_s),
        .c_out(fa_s3_c57_n76_c)
    );

    fa fa_s3_c57_n77 (
        .a(stage3_col57[6]),
        .b(stage3_col57[7]),
        .c_in(stage3_col57[8]),
        .s(fa_s3_c57_n77_s),
        .c_out(fa_s3_c57_n77_c)
    );

    fa fa_s3_c58_n78 (
        .a(stage3_col58[0]),
        .b(stage3_col58[1]),
        .c_in(stage3_col58[2]),
        .s(fa_s3_c58_n78_s),
        .c_out(fa_s3_c58_n78_c)
    );

    fa fa_s3_c58_n79 (
        .a(stage3_col58[3]),
        .b(stage3_col58[4]),
        .c_in(stage3_col58[5]),
        .s(fa_s3_c58_n79_s),
        .c_out(fa_s3_c58_n79_c)
    );

    fa fa_s3_c58_n80 (
        .a(stage3_col58[6]),
        .b(stage3_col58[7]),
        .c_in(stage3_col58[8]),
        .s(fa_s3_c58_n80_s),
        .c_out(fa_s3_c58_n80_c)
    );

    fa fa_s3_c59_n81 (
        .a(stage3_col59[0]),
        .b(stage3_col59[1]),
        .c_in(stage3_col59[2]),
        .s(fa_s3_c59_n81_s),
        .c_out(fa_s3_c59_n81_c)
    );

    fa fa_s3_c59_n82 (
        .a(stage3_col59[3]),
        .b(stage3_col59[4]),
        .c_in(stage3_col59[5]),
        .s(fa_s3_c59_n82_s),
        .c_out(fa_s3_c59_n82_c)
    );

    fa fa_s3_c59_n83 (
        .a(stage3_col59[6]),
        .b(stage3_col59[7]),
        .c_in(stage3_col59[8]),
        .s(fa_s3_c59_n83_s),
        .c_out(fa_s3_c59_n83_c)
    );

    fa fa_s3_c60_n84 (
        .a(stage3_col60[0]),
        .b(stage3_col60[1]),
        .c_in(stage3_col60[2]),
        .s(fa_s3_c60_n84_s),
        .c_out(fa_s3_c60_n84_c)
    );

    fa fa_s3_c60_n85 (
        .a(stage3_col60[3]),
        .b(stage3_col60[4]),
        .c_in(stage3_col60[5]),
        .s(fa_s3_c60_n85_s),
        .c_out(fa_s3_c60_n85_c)
    );

    fa fa_s3_c60_n86 (
        .a(stage3_col60[6]),
        .b(stage3_col60[7]),
        .c_in(stage3_col60[8]),
        .s(fa_s3_c60_n86_s),
        .c_out(fa_s3_c60_n86_c)
    );

    fa fa_s3_c61_n87 (
        .a(stage3_col61[0]),
        .b(stage3_col61[1]),
        .c_in(stage3_col61[2]),
        .s(fa_s3_c61_n87_s),
        .c_out(fa_s3_c61_n87_c)
    );

    fa fa_s3_c61_n88 (
        .a(stage3_col61[3]),
        .b(stage3_col61[4]),
        .c_in(stage3_col61[5]),
        .s(fa_s3_c61_n88_s),
        .c_out(fa_s3_c61_n88_c)
    );

    fa fa_s3_c61_n89 (
        .a(stage3_col61[6]),
        .b(stage3_col61[7]),
        .c_in(stage3_col61[8]),
        .s(fa_s3_c61_n89_s),
        .c_out(fa_s3_c61_n89_c)
    );

    fa fa_s3_c62_n90 (
        .a(stage3_col62[0]),
        .b(stage3_col62[1]),
        .c_in(stage3_col62[2]),
        .s(fa_s3_c62_n90_s),
        .c_out(fa_s3_c62_n90_c)
    );

    fa fa_s3_c62_n91 (
        .a(stage3_col62[3]),
        .b(stage3_col62[4]),
        .c_in(stage3_col62[5]),
        .s(fa_s3_c62_n91_s),
        .c_out(fa_s3_c62_n91_c)
    );

    fa fa_s3_c62_n92 (
        .a(stage3_col62[6]),
        .b(stage3_col62[7]),
        .c_in(stage3_col62[8]),
        .s(fa_s3_c62_n92_s),
        .c_out(fa_s3_c62_n92_c)
    );

    fa fa_s3_c63_n93 (
        .a(stage3_col63[0]),
        .b(stage3_col63[1]),
        .c_in(stage3_col63[2]),
        .s(fa_s3_c63_n93_s),
        .c_out(fa_s3_c63_n93_c)
    );

    fa fa_s3_c63_n94 (
        .a(stage3_col63[3]),
        .b(stage3_col63[4]),
        .c_in(stage3_col63[5]),
        .s(fa_s3_c63_n94_s),
        .c_out(fa_s3_c63_n94_c)
    );

    fa fa_s3_c63_n95 (
        .a(stage3_col63[6]),
        .b(stage3_col63[7]),
        .c_in(stage3_col63[8]),
        .s(fa_s3_c63_n95_s),
        .c_out(fa_s3_c63_n95_c)
    );

    fa fa_s3_c64_n96 (
        .a(stage3_col64[0]),
        .b(stage3_col64[1]),
        .c_in(stage3_col64[2]),
        .s(fa_s3_c64_n96_s),
        .c_out(fa_s3_c64_n96_c)
    );

    fa fa_s3_c64_n97 (
        .a(stage3_col64[3]),
        .b(stage3_col64[4]),
        .c_in(stage3_col64[5]),
        .s(fa_s3_c64_n97_s),
        .c_out(fa_s3_c64_n97_c)
    );

    fa fa_s3_c64_n98 (
        .a(stage3_col64[6]),
        .b(stage3_col64[7]),
        .c_in(stage3_col64[8]),
        .s(fa_s3_c64_n98_s),
        .c_out(fa_s3_c64_n98_c)
    );

    fa fa_s3_c65_n99 (
        .a(stage3_col65[0]),
        .b(stage3_col65[1]),
        .c_in(stage3_col65[2]),
        .s(fa_s3_c65_n99_s),
        .c_out(fa_s3_c65_n99_c)
    );

    fa fa_s3_c65_n100 (
        .a(stage3_col65[3]),
        .b(stage3_col65[4]),
        .c_in(stage3_col65[5]),
        .s(fa_s3_c65_n100_s),
        .c_out(fa_s3_c65_n100_c)
    );

    fa fa_s3_c65_n101 (
        .a(stage3_col65[6]),
        .b(stage3_col65[7]),
        .c_in(stage3_col65[8]),
        .s(fa_s3_c65_n101_s),
        .c_out(fa_s3_c65_n101_c)
    );

    fa fa_s3_c66_n102 (
        .a(stage3_col66[0]),
        .b(stage3_col66[1]),
        .c_in(stage3_col66[2]),
        .s(fa_s3_c66_n102_s),
        .c_out(fa_s3_c66_n102_c)
    );

    fa fa_s3_c66_n103 (
        .a(stage3_col66[3]),
        .b(stage3_col66[4]),
        .c_in(stage3_col66[5]),
        .s(fa_s3_c66_n103_s),
        .c_out(fa_s3_c66_n103_c)
    );

    fa fa_s3_c66_n104 (
        .a(stage3_col66[6]),
        .b(stage3_col66[7]),
        .c_in(stage3_col66[8]),
        .s(fa_s3_c66_n104_s),
        .c_out(fa_s3_c66_n104_c)
    );

    fa fa_s3_c67_n105 (
        .a(stage3_col67[0]),
        .b(stage3_col67[1]),
        .c_in(stage3_col67[2]),
        .s(fa_s3_c67_n105_s),
        .c_out(fa_s3_c67_n105_c)
    );

    fa fa_s3_c67_n106 (
        .a(stage3_col67[3]),
        .b(stage3_col67[4]),
        .c_in(stage3_col67[5]),
        .s(fa_s3_c67_n106_s),
        .c_out(fa_s3_c67_n106_c)
    );

    fa fa_s3_c67_n107 (
        .a(stage3_col67[6]),
        .b(stage3_col67[7]),
        .c_in(stage3_col67[8]),
        .s(fa_s3_c67_n107_s),
        .c_out(fa_s3_c67_n107_c)
    );

    fa fa_s3_c68_n108 (
        .a(stage3_col68[0]),
        .b(stage3_col68[1]),
        .c_in(stage3_col68[2]),
        .s(fa_s3_c68_n108_s),
        .c_out(fa_s3_c68_n108_c)
    );

    fa fa_s3_c68_n109 (
        .a(stage3_col68[3]),
        .b(stage3_col68[4]),
        .c_in(stage3_col68[5]),
        .s(fa_s3_c68_n109_s),
        .c_out(fa_s3_c68_n109_c)
    );

    fa fa_s3_c68_n110 (
        .a(stage3_col68[6]),
        .b(stage3_col68[7]),
        .c_in(stage3_col68[8]),
        .s(fa_s3_c68_n110_s),
        .c_out(fa_s3_c68_n110_c)
    );

    fa fa_s3_c69_n111 (
        .a(stage3_col69[0]),
        .b(stage3_col69[1]),
        .c_in(stage3_col69[2]),
        .s(fa_s3_c69_n111_s),
        .c_out(fa_s3_c69_n111_c)
    );

    fa fa_s3_c69_n112 (
        .a(stage3_col69[3]),
        .b(stage3_col69[4]),
        .c_in(stage3_col69[5]),
        .s(fa_s3_c69_n112_s),
        .c_out(fa_s3_c69_n112_c)
    );

    fa fa_s3_c69_n113 (
        .a(stage3_col69[6]),
        .b(stage3_col69[7]),
        .c_in(stage3_col69[8]),
        .s(fa_s3_c69_n113_s),
        .c_out(fa_s3_c69_n113_c)
    );

    fa fa_s3_c70_n114 (
        .a(stage3_col70[0]),
        .b(stage3_col70[1]),
        .c_in(stage3_col70[2]),
        .s(fa_s3_c70_n114_s),
        .c_out(fa_s3_c70_n114_c)
    );

    fa fa_s3_c70_n115 (
        .a(stage3_col70[3]),
        .b(stage3_col70[4]),
        .c_in(stage3_col70[5]),
        .s(fa_s3_c70_n115_s),
        .c_out(fa_s3_c70_n115_c)
    );

    fa fa_s3_c70_n116 (
        .a(stage3_col70[6]),
        .b(stage3_col70[7]),
        .c_in(stage3_col70[8]),
        .s(fa_s3_c70_n116_s),
        .c_out(fa_s3_c70_n116_c)
    );

    fa fa_s3_c71_n117 (
        .a(stage3_col71[0]),
        .b(stage3_col71[1]),
        .c_in(stage3_col71[2]),
        .s(fa_s3_c71_n117_s),
        .c_out(fa_s3_c71_n117_c)
    );

    fa fa_s3_c71_n118 (
        .a(stage3_col71[3]),
        .b(stage3_col71[4]),
        .c_in(stage3_col71[5]),
        .s(fa_s3_c71_n118_s),
        .c_out(fa_s3_c71_n118_c)
    );

    fa fa_s3_c71_n119 (
        .a(stage3_col71[6]),
        .b(stage3_col71[7]),
        .c_in(stage3_col71[8]),
        .s(fa_s3_c71_n119_s),
        .c_out(fa_s3_c71_n119_c)
    );

    fa fa_s3_c72_n120 (
        .a(stage3_col72[0]),
        .b(stage3_col72[1]),
        .c_in(stage3_col72[2]),
        .s(fa_s3_c72_n120_s),
        .c_out(fa_s3_c72_n120_c)
    );

    fa fa_s3_c72_n121 (
        .a(stage3_col72[3]),
        .b(stage3_col72[4]),
        .c_in(stage3_col72[5]),
        .s(fa_s3_c72_n121_s),
        .c_out(fa_s3_c72_n121_c)
    );

    fa fa_s3_c72_n122 (
        .a(stage3_col72[6]),
        .b(stage3_col72[7]),
        .c_in(stage3_col72[8]),
        .s(fa_s3_c72_n122_s),
        .c_out(fa_s3_c72_n122_c)
    );

    fa fa_s3_c73_n123 (
        .a(stage3_col73[0]),
        .b(stage3_col73[1]),
        .c_in(stage3_col73[2]),
        .s(fa_s3_c73_n123_s),
        .c_out(fa_s3_c73_n123_c)
    );

    fa fa_s3_c73_n124 (
        .a(stage3_col73[3]),
        .b(stage3_col73[4]),
        .c_in(stage3_col73[5]),
        .s(fa_s3_c73_n124_s),
        .c_out(fa_s3_c73_n124_c)
    );

    fa fa_s3_c73_n125 (
        .a(stage3_col73[6]),
        .b(stage3_col73[7]),
        .c_in(stage3_col73[8]),
        .s(fa_s3_c73_n125_s),
        .c_out(fa_s3_c73_n125_c)
    );

    fa fa_s3_c74_n126 (
        .a(stage3_col74[0]),
        .b(stage3_col74[1]),
        .c_in(stage3_col74[2]),
        .s(fa_s3_c74_n126_s),
        .c_out(fa_s3_c74_n126_c)
    );

    fa fa_s3_c74_n127 (
        .a(stage3_col74[3]),
        .b(stage3_col74[4]),
        .c_in(stage3_col74[5]),
        .s(fa_s3_c74_n127_s),
        .c_out(fa_s3_c74_n127_c)
    );

    fa fa_s3_c74_n128 (
        .a(stage3_col74[6]),
        .b(stage3_col74[7]),
        .c_in(stage3_col74[8]),
        .s(fa_s3_c74_n128_s),
        .c_out(fa_s3_c74_n128_c)
    );

    fa fa_s3_c75_n129 (
        .a(stage3_col75[0]),
        .b(stage3_col75[1]),
        .c_in(stage3_col75[2]),
        .s(fa_s3_c75_n129_s),
        .c_out(fa_s3_c75_n129_c)
    );

    fa fa_s3_c75_n130 (
        .a(stage3_col75[3]),
        .b(stage3_col75[4]),
        .c_in(stage3_col75[5]),
        .s(fa_s3_c75_n130_s),
        .c_out(fa_s3_c75_n130_c)
    );

    fa fa_s3_c75_n131 (
        .a(stage3_col75[6]),
        .b(stage3_col75[7]),
        .c_in(stage3_col75[8]),
        .s(fa_s3_c75_n131_s),
        .c_out(fa_s3_c75_n131_c)
    );

    fa fa_s3_c76_n132 (
        .a(stage3_col76[0]),
        .b(stage3_col76[1]),
        .c_in(stage3_col76[2]),
        .s(fa_s3_c76_n132_s),
        .c_out(fa_s3_c76_n132_c)
    );

    fa fa_s3_c76_n133 (
        .a(stage3_col76[3]),
        .b(stage3_col76[4]),
        .c_in(stage3_col76[5]),
        .s(fa_s3_c76_n133_s),
        .c_out(fa_s3_c76_n133_c)
    );

    fa fa_s3_c76_n134 (
        .a(stage3_col76[6]),
        .b(stage3_col76[7]),
        .c_in(stage3_col76[8]),
        .s(fa_s3_c76_n134_s),
        .c_out(fa_s3_c76_n134_c)
    );

    fa fa_s3_c77_n135 (
        .a(stage3_col77[0]),
        .b(stage3_col77[1]),
        .c_in(stage3_col77[2]),
        .s(fa_s3_c77_n135_s),
        .c_out(fa_s3_c77_n135_c)
    );

    fa fa_s3_c77_n136 (
        .a(stage3_col77[3]),
        .b(stage3_col77[4]),
        .c_in(stage3_col77[5]),
        .s(fa_s3_c77_n136_s),
        .c_out(fa_s3_c77_n136_c)
    );

    fa fa_s3_c77_n137 (
        .a(stage3_col77[6]),
        .b(stage3_col77[7]),
        .c_in(stage3_col77[8]),
        .s(fa_s3_c77_n137_s),
        .c_out(fa_s3_c77_n137_c)
    );

    fa fa_s3_c78_n138 (
        .a(stage3_col78[0]),
        .b(stage3_col78[1]),
        .c_in(stage3_col78[2]),
        .s(fa_s3_c78_n138_s),
        .c_out(fa_s3_c78_n138_c)
    );

    fa fa_s3_c78_n139 (
        .a(stage3_col78[3]),
        .b(stage3_col78[4]),
        .c_in(stage3_col78[5]),
        .s(fa_s3_c78_n139_s),
        .c_out(fa_s3_c78_n139_c)
    );

    fa fa_s3_c78_n140 (
        .a(stage3_col78[6]),
        .b(stage3_col78[7]),
        .c_in(stage3_col78[8]),
        .s(fa_s3_c78_n140_s),
        .c_out(fa_s3_c78_n140_c)
    );

    fa fa_s3_c79_n141 (
        .a(stage3_col79[0]),
        .b(stage3_col79[1]),
        .c_in(stage3_col79[2]),
        .s(fa_s3_c79_n141_s),
        .c_out(fa_s3_c79_n141_c)
    );

    fa fa_s3_c79_n142 (
        .a(stage3_col79[3]),
        .b(stage3_col79[4]),
        .c_in(stage3_col79[5]),
        .s(fa_s3_c79_n142_s),
        .c_out(fa_s3_c79_n142_c)
    );

    fa fa_s3_c79_n143 (
        .a(stage3_col79[6]),
        .b(stage3_col79[7]),
        .c_in(stage3_col79[8]),
        .s(fa_s3_c79_n143_s),
        .c_out(fa_s3_c79_n143_c)
    );

    fa fa_s3_c80_n144 (
        .a(stage3_col80[0]),
        .b(stage3_col80[1]),
        .c_in(stage3_col80[2]),
        .s(fa_s3_c80_n144_s),
        .c_out(fa_s3_c80_n144_c)
    );

    fa fa_s3_c80_n145 (
        .a(stage3_col80[3]),
        .b(stage3_col80[4]),
        .c_in(stage3_col80[5]),
        .s(fa_s3_c80_n145_s),
        .c_out(fa_s3_c80_n145_c)
    );

    fa fa_s3_c80_n146 (
        .a(stage3_col80[6]),
        .b(stage3_col80[7]),
        .c_in(stage3_col80[8]),
        .s(fa_s3_c80_n146_s),
        .c_out(fa_s3_c80_n146_c)
    );

    fa fa_s3_c81_n147 (
        .a(stage3_col81[0]),
        .b(stage3_col81[1]),
        .c_in(stage3_col81[2]),
        .s(fa_s3_c81_n147_s),
        .c_out(fa_s3_c81_n147_c)
    );

    fa fa_s3_c81_n148 (
        .a(stage3_col81[3]),
        .b(stage3_col81[4]),
        .c_in(stage3_col81[5]),
        .s(fa_s3_c81_n148_s),
        .c_out(fa_s3_c81_n148_c)
    );

    fa fa_s3_c81_n149 (
        .a(stage3_col81[6]),
        .b(stage3_col81[7]),
        .c_in(stage3_col81[8]),
        .s(fa_s3_c81_n149_s),
        .c_out(fa_s3_c81_n149_c)
    );

    fa fa_s3_c82_n150 (
        .a(stage3_col82[0]),
        .b(stage3_col82[1]),
        .c_in(stage3_col82[2]),
        .s(fa_s3_c82_n150_s),
        .c_out(fa_s3_c82_n150_c)
    );

    fa fa_s3_c82_n151 (
        .a(stage3_col82[3]),
        .b(stage3_col82[4]),
        .c_in(stage3_col82[5]),
        .s(fa_s3_c82_n151_s),
        .c_out(fa_s3_c82_n151_c)
    );

    fa fa_s3_c82_n152 (
        .a(stage3_col82[6]),
        .b(stage3_col82[7]),
        .c_in(stage3_col82[8]),
        .s(fa_s3_c82_n152_s),
        .c_out(fa_s3_c82_n152_c)
    );

    fa fa_s3_c83_n153 (
        .a(stage3_col83[0]),
        .b(stage3_col83[1]),
        .c_in(stage3_col83[2]),
        .s(fa_s3_c83_n153_s),
        .c_out(fa_s3_c83_n153_c)
    );

    fa fa_s3_c83_n154 (
        .a(stage3_col83[3]),
        .b(stage3_col83[4]),
        .c_in(stage3_col83[5]),
        .s(fa_s3_c83_n154_s),
        .c_out(fa_s3_c83_n154_c)
    );

    fa fa_s3_c83_n155 (
        .a(stage3_col83[6]),
        .b(stage3_col83[7]),
        .c_in(stage3_col83[8]),
        .s(fa_s3_c83_n155_s),
        .c_out(fa_s3_c83_n155_c)
    );

    fa fa_s3_c84_n156 (
        .a(stage3_col84[0]),
        .b(stage3_col84[1]),
        .c_in(stage3_col84[2]),
        .s(fa_s3_c84_n156_s),
        .c_out(fa_s3_c84_n156_c)
    );

    fa fa_s3_c84_n157 (
        .a(stage3_col84[3]),
        .b(stage3_col84[4]),
        .c_in(stage3_col84[5]),
        .s(fa_s3_c84_n157_s),
        .c_out(fa_s3_c84_n157_c)
    );

    fa fa_s3_c84_n158 (
        .a(stage3_col84[6]),
        .b(stage3_col84[7]),
        .c_in(stage3_col84[8]),
        .s(fa_s3_c84_n158_s),
        .c_out(fa_s3_c84_n158_c)
    );

    fa fa_s3_c85_n159 (
        .a(stage3_col85[0]),
        .b(stage3_col85[1]),
        .c_in(stage3_col85[2]),
        .s(fa_s3_c85_n159_s),
        .c_out(fa_s3_c85_n159_c)
    );

    fa fa_s3_c85_n160 (
        .a(stage3_col85[3]),
        .b(stage3_col85[4]),
        .c_in(stage3_col85[5]),
        .s(fa_s3_c85_n160_s),
        .c_out(fa_s3_c85_n160_c)
    );

    fa fa_s3_c85_n161 (
        .a(stage3_col85[6]),
        .b(stage3_col85[7]),
        .c_in(stage3_col85[8]),
        .s(fa_s3_c85_n161_s),
        .c_out(fa_s3_c85_n161_c)
    );

    fa fa_s3_c86_n162 (
        .a(stage3_col86[0]),
        .b(stage3_col86[1]),
        .c_in(stage3_col86[2]),
        .s(fa_s3_c86_n162_s),
        .c_out(fa_s3_c86_n162_c)
    );

    fa fa_s3_c86_n163 (
        .a(stage3_col86[3]),
        .b(stage3_col86[4]),
        .c_in(stage3_col86[5]),
        .s(fa_s3_c86_n163_s),
        .c_out(fa_s3_c86_n163_c)
    );

    fa fa_s3_c86_n164 (
        .a(stage3_col86[6]),
        .b(stage3_col86[7]),
        .c_in(stage3_col86[8]),
        .s(fa_s3_c86_n164_s),
        .c_out(fa_s3_c86_n164_c)
    );

    fa fa_s3_c87_n165 (
        .a(stage3_col87[0]),
        .b(stage3_col87[1]),
        .c_in(stage3_col87[2]),
        .s(fa_s3_c87_n165_s),
        .c_out(fa_s3_c87_n165_c)
    );

    fa fa_s3_c87_n166 (
        .a(stage3_col87[3]),
        .b(stage3_col87[4]),
        .c_in(stage3_col87[5]),
        .s(fa_s3_c87_n166_s),
        .c_out(fa_s3_c87_n166_c)
    );

    fa fa_s3_c87_n167 (
        .a(stage3_col87[6]),
        .b(stage3_col87[7]),
        .c_in(stage3_col87[8]),
        .s(fa_s3_c87_n167_s),
        .c_out(fa_s3_c87_n167_c)
    );

    fa fa_s3_c88_n168 (
        .a(stage3_col88[0]),
        .b(stage3_col88[1]),
        .c_in(stage3_col88[2]),
        .s(fa_s3_c88_n168_s),
        .c_out(fa_s3_c88_n168_c)
    );

    fa fa_s3_c88_n169 (
        .a(stage3_col88[3]),
        .b(stage3_col88[4]),
        .c_in(stage3_col88[5]),
        .s(fa_s3_c88_n169_s),
        .c_out(fa_s3_c88_n169_c)
    );

    fa fa_s3_c88_n170 (
        .a(stage3_col88[6]),
        .b(stage3_col88[7]),
        .c_in(stage3_col88[8]),
        .s(fa_s3_c88_n170_s),
        .c_out(fa_s3_c88_n170_c)
    );

    fa fa_s3_c89_n171 (
        .a(stage3_col89[0]),
        .b(stage3_col89[1]),
        .c_in(stage3_col89[2]),
        .s(fa_s3_c89_n171_s),
        .c_out(fa_s3_c89_n171_c)
    );

    fa fa_s3_c89_n172 (
        .a(stage3_col89[3]),
        .b(stage3_col89[4]),
        .c_in(stage3_col89[5]),
        .s(fa_s3_c89_n172_s),
        .c_out(fa_s3_c89_n172_c)
    );

    fa fa_s3_c89_n173 (
        .a(stage3_col89[6]),
        .b(stage3_col89[7]),
        .c_in(stage3_col89[8]),
        .s(fa_s3_c89_n173_s),
        .c_out(fa_s3_c89_n173_c)
    );

    fa fa_s3_c90_n174 (
        .a(stage3_col90[0]),
        .b(stage3_col90[1]),
        .c_in(stage3_col90[2]),
        .s(fa_s3_c90_n174_s),
        .c_out(fa_s3_c90_n174_c)
    );

    fa fa_s3_c90_n175 (
        .a(stage3_col90[3]),
        .b(stage3_col90[4]),
        .c_in(stage3_col90[5]),
        .s(fa_s3_c90_n175_s),
        .c_out(fa_s3_c90_n175_c)
    );

    fa fa_s3_c90_n176 (
        .a(stage3_col90[6]),
        .b(stage3_col90[7]),
        .c_in(stage3_col90[8]),
        .s(fa_s3_c90_n176_s),
        .c_out(fa_s3_c90_n176_c)
    );

    fa fa_s3_c91_n177 (
        .a(stage3_col91[0]),
        .b(stage3_col91[1]),
        .c_in(stage3_col91[2]),
        .s(fa_s3_c91_n177_s),
        .c_out(fa_s3_c91_n177_c)
    );

    fa fa_s3_c91_n178 (
        .a(stage3_col91[3]),
        .b(stage3_col91[4]),
        .c_in(stage3_col91[5]),
        .s(fa_s3_c91_n178_s),
        .c_out(fa_s3_c91_n178_c)
    );

    fa fa_s3_c91_n179 (
        .a(stage3_col91[6]),
        .b(stage3_col91[7]),
        .c_in(stage3_col91[8]),
        .s(fa_s3_c91_n179_s),
        .c_out(fa_s3_c91_n179_c)
    );

    fa fa_s3_c92_n180 (
        .a(stage3_col92[0]),
        .b(stage3_col92[1]),
        .c_in(stage3_col92[2]),
        .s(fa_s3_c92_n180_s),
        .c_out(fa_s3_c92_n180_c)
    );

    fa fa_s3_c92_n181 (
        .a(stage3_col92[3]),
        .b(stage3_col92[4]),
        .c_in(stage3_col92[5]),
        .s(fa_s3_c92_n181_s),
        .c_out(fa_s3_c92_n181_c)
    );

    fa fa_s3_c92_n182 (
        .a(stage3_col92[6]),
        .b(stage3_col92[7]),
        .c_in(stage3_col92[8]),
        .s(fa_s3_c92_n182_s),
        .c_out(fa_s3_c92_n182_c)
    );

    fa fa_s3_c93_n183 (
        .a(stage3_col93[0]),
        .b(stage3_col93[1]),
        .c_in(stage3_col93[2]),
        .s(fa_s3_c93_n183_s),
        .c_out(fa_s3_c93_n183_c)
    );

    fa fa_s3_c93_n184 (
        .a(stage3_col93[3]),
        .b(stage3_col93[4]),
        .c_in(stage3_col93[5]),
        .s(fa_s3_c93_n184_s),
        .c_out(fa_s3_c93_n184_c)
    );

    fa fa_s3_c93_n185 (
        .a(stage3_col93[6]),
        .b(stage3_col93[7]),
        .c_in(stage3_col93[8]),
        .s(fa_s3_c93_n185_s),
        .c_out(fa_s3_c93_n185_c)
    );

    fa fa_s3_c94_n186 (
        .a(stage3_col94[0]),
        .b(stage3_col94[1]),
        .c_in(stage3_col94[2]),
        .s(fa_s3_c94_n186_s),
        .c_out(fa_s3_c94_n186_c)
    );

    fa fa_s3_c94_n187 (
        .a(stage3_col94[3]),
        .b(stage3_col94[4]),
        .c_in(stage3_col94[5]),
        .s(fa_s3_c94_n187_s),
        .c_out(fa_s3_c94_n187_c)
    );

    fa fa_s3_c94_n188 (
        .a(stage3_col94[6]),
        .b(stage3_col94[7]),
        .c_in(stage3_col94[8]),
        .s(fa_s3_c94_n188_s),
        .c_out(fa_s3_c94_n188_c)
    );

    fa fa_s3_c95_n189 (
        .a(stage3_col95[0]),
        .b(stage3_col95[1]),
        .c_in(stage3_col95[2]),
        .s(fa_s3_c95_n189_s),
        .c_out(fa_s3_c95_n189_c)
    );

    fa fa_s3_c95_n190 (
        .a(stage3_col95[3]),
        .b(stage3_col95[4]),
        .c_in(stage3_col95[5]),
        .s(fa_s3_c95_n190_s),
        .c_out(fa_s3_c95_n190_c)
    );

    fa fa_s3_c95_n191 (
        .a(stage3_col95[6]),
        .b(stage3_col95[7]),
        .c_in(stage3_col95[8]),
        .s(fa_s3_c95_n191_s),
        .c_out(fa_s3_c95_n191_c)
    );

    fa fa_s3_c96_n192 (
        .a(stage3_col96[0]),
        .b(stage3_col96[1]),
        .c_in(stage3_col96[2]),
        .s(fa_s3_c96_n192_s),
        .c_out(fa_s3_c96_n192_c)
    );

    fa fa_s3_c96_n193 (
        .a(stage3_col96[3]),
        .b(stage3_col96[4]),
        .c_in(stage3_col96[5]),
        .s(fa_s3_c96_n193_s),
        .c_out(fa_s3_c96_n193_c)
    );

    fa fa_s3_c96_n194 (
        .a(stage3_col96[6]),
        .b(stage3_col96[7]),
        .c_in(stage3_col96[8]),
        .s(fa_s3_c96_n194_s),
        .c_out(fa_s3_c96_n194_c)
    );

    fa fa_s3_c97_n195 (
        .a(stage3_col97[0]),
        .b(stage3_col97[1]),
        .c_in(stage3_col97[2]),
        .s(fa_s3_c97_n195_s),
        .c_out(fa_s3_c97_n195_c)
    );

    fa fa_s3_c97_n196 (
        .a(stage3_col97[3]),
        .b(stage3_col97[4]),
        .c_in(stage3_col97[5]),
        .s(fa_s3_c97_n196_s),
        .c_out(fa_s3_c97_n196_c)
    );

    fa fa_s3_c97_n197 (
        .a(stage3_col97[6]),
        .b(stage3_col97[7]),
        .c_in(stage3_col97[8]),
        .s(fa_s3_c97_n197_s),
        .c_out(fa_s3_c97_n197_c)
    );

    fa fa_s3_c98_n198 (
        .a(stage3_col98[0]),
        .b(stage3_col98[1]),
        .c_in(stage3_col98[2]),
        .s(fa_s3_c98_n198_s),
        .c_out(fa_s3_c98_n198_c)
    );

    fa fa_s3_c98_n199 (
        .a(stage3_col98[3]),
        .b(stage3_col98[4]),
        .c_in(stage3_col98[5]),
        .s(fa_s3_c98_n199_s),
        .c_out(fa_s3_c98_n199_c)
    );

    fa fa_s3_c98_n200 (
        .a(stage3_col98[6]),
        .b(stage3_col98[7]),
        .c_in(stage3_col98[8]),
        .s(fa_s3_c98_n200_s),
        .c_out(fa_s3_c98_n200_c)
    );

    fa fa_s3_c99_n201 (
        .a(stage3_col99[0]),
        .b(stage3_col99[1]),
        .c_in(stage3_col99[2]),
        .s(fa_s3_c99_n201_s),
        .c_out(fa_s3_c99_n201_c)
    );

    fa fa_s3_c99_n202 (
        .a(stage3_col99[3]),
        .b(stage3_col99[4]),
        .c_in(stage3_col99[5]),
        .s(fa_s3_c99_n202_s),
        .c_out(fa_s3_c99_n202_c)
    );

    fa fa_s3_c99_n203 (
        .a(stage3_col99[6]),
        .b(stage3_col99[7]),
        .c_in(stage3_col99[8]),
        .s(fa_s3_c99_n203_s),
        .c_out(fa_s3_c99_n203_c)
    );

    fa fa_s3_c100_n204 (
        .a(stage3_col100[0]),
        .b(stage3_col100[1]),
        .c_in(stage3_col100[2]),
        .s(fa_s3_c100_n204_s),
        .c_out(fa_s3_c100_n204_c)
    );

    fa fa_s3_c100_n205 (
        .a(stage3_col100[3]),
        .b(stage3_col100[4]),
        .c_in(stage3_col100[5]),
        .s(fa_s3_c100_n205_s),
        .c_out(fa_s3_c100_n205_c)
    );

    fa fa_s3_c100_n206 (
        .a(stage3_col100[6]),
        .b(stage3_col100[7]),
        .c_in(stage3_col100[8]),
        .s(fa_s3_c100_n206_s),
        .c_out(fa_s3_c100_n206_c)
    );

    fa fa_s3_c101_n207 (
        .a(stage3_col101[0]),
        .b(stage3_col101[1]),
        .c_in(stage3_col101[2]),
        .s(fa_s3_c101_n207_s),
        .c_out(fa_s3_c101_n207_c)
    );

    fa fa_s3_c101_n208 (
        .a(stage3_col101[3]),
        .b(stage3_col101[4]),
        .c_in(stage3_col101[5]),
        .s(fa_s3_c101_n208_s),
        .c_out(fa_s3_c101_n208_c)
    );

    fa fa_s3_c101_n209 (
        .a(stage3_col101[6]),
        .b(stage3_col101[7]),
        .c_in(stage3_col101[8]),
        .s(fa_s3_c101_n209_s),
        .c_out(fa_s3_c101_n209_c)
    );

    fa fa_s3_c102_n210 (
        .a(stage3_col102[0]),
        .b(stage3_col102[1]),
        .c_in(stage3_col102[2]),
        .s(fa_s3_c102_n210_s),
        .c_out(fa_s3_c102_n210_c)
    );

    fa fa_s3_c102_n211 (
        .a(stage3_col102[3]),
        .b(stage3_col102[4]),
        .c_in(stage3_col102[5]),
        .s(fa_s3_c102_n211_s),
        .c_out(fa_s3_c102_n211_c)
    );

    fa fa_s3_c102_n212 (
        .a(stage3_col102[6]),
        .b(stage3_col102[7]),
        .c_in(stage3_col102[8]),
        .s(fa_s3_c102_n212_s),
        .c_out(fa_s3_c102_n212_c)
    );

    fa fa_s3_c103_n213 (
        .a(stage3_col103[0]),
        .b(stage3_col103[1]),
        .c_in(stage3_col103[2]),
        .s(fa_s3_c103_n213_s),
        .c_out(fa_s3_c103_n213_c)
    );

    fa fa_s3_c103_n214 (
        .a(stage3_col103[3]),
        .b(stage3_col103[4]),
        .c_in(stage3_col103[5]),
        .s(fa_s3_c103_n214_s),
        .c_out(fa_s3_c103_n214_c)
    );

    fa fa_s3_c103_n215 (
        .a(stage3_col103[6]),
        .b(stage3_col103[7]),
        .c_in(stage3_col103[8]),
        .s(fa_s3_c103_n215_s),
        .c_out(fa_s3_c103_n215_c)
    );

    fa fa_s3_c104_n216 (
        .a(stage3_col104[0]),
        .b(stage3_col104[1]),
        .c_in(stage3_col104[2]),
        .s(fa_s3_c104_n216_s),
        .c_out(fa_s3_c104_n216_c)
    );

    fa fa_s3_c104_n217 (
        .a(stage3_col104[3]),
        .b(stage3_col104[4]),
        .c_in(stage3_col104[5]),
        .s(fa_s3_c104_n217_s),
        .c_out(fa_s3_c104_n217_c)
    );

    fa fa_s3_c104_n218 (
        .a(stage3_col104[6]),
        .b(stage3_col104[7]),
        .c_in(stage3_col104[8]),
        .s(fa_s3_c104_n218_s),
        .c_out(fa_s3_c104_n218_c)
    );

    fa fa_s3_c105_n219 (
        .a(stage3_col105[0]),
        .b(stage3_col105[1]),
        .c_in(stage3_col105[2]),
        .s(fa_s3_c105_n219_s),
        .c_out(fa_s3_c105_n219_c)
    );

    fa fa_s3_c105_n220 (
        .a(stage3_col105[3]),
        .b(stage3_col105[4]),
        .c_in(stage3_col105[5]),
        .s(fa_s3_c105_n220_s),
        .c_out(fa_s3_c105_n220_c)
    );

    fa fa_s3_c105_n221 (
        .a(stage3_col105[6]),
        .b(stage3_col105[7]),
        .c_in(stage3_col105[8]),
        .s(fa_s3_c105_n221_s),
        .c_out(fa_s3_c105_n221_c)
    );

    fa fa_s3_c106_n222 (
        .a(stage3_col106[0]),
        .b(stage3_col106[1]),
        .c_in(stage3_col106[2]),
        .s(fa_s3_c106_n222_s),
        .c_out(fa_s3_c106_n222_c)
    );

    fa fa_s3_c106_n223 (
        .a(stage3_col106[3]),
        .b(stage3_col106[4]),
        .c_in(stage3_col106[5]),
        .s(fa_s3_c106_n223_s),
        .c_out(fa_s3_c106_n223_c)
    );

    fa fa_s3_c106_n224 (
        .a(stage3_col106[6]),
        .b(stage3_col106[7]),
        .c_in(stage3_col106[8]),
        .s(fa_s3_c106_n224_s),
        .c_out(fa_s3_c106_n224_c)
    );

    fa fa_s3_c107_n225 (
        .a(stage3_col107[0]),
        .b(stage3_col107[1]),
        .c_in(stage3_col107[2]),
        .s(fa_s3_c107_n225_s),
        .c_out(fa_s3_c107_n225_c)
    );

    fa fa_s3_c107_n226 (
        .a(stage3_col107[3]),
        .b(stage3_col107[4]),
        .c_in(stage3_col107[5]),
        .s(fa_s3_c107_n226_s),
        .c_out(fa_s3_c107_n226_c)
    );

    fa fa_s3_c107_n227 (
        .a(stage3_col107[6]),
        .b(stage3_col107[7]),
        .c_in(stage3_col107[8]),
        .s(fa_s3_c107_n227_s),
        .c_out(fa_s3_c107_n227_c)
    );

    fa fa_s3_c108_n228 (
        .a(stage3_col108[0]),
        .b(stage3_col108[1]),
        .c_in(stage3_col108[2]),
        .s(fa_s3_c108_n228_s),
        .c_out(fa_s3_c108_n228_c)
    );

    fa fa_s3_c108_n229 (
        .a(stage3_col108[3]),
        .b(stage3_col108[4]),
        .c_in(stage3_col108[5]),
        .s(fa_s3_c108_n229_s),
        .c_out(fa_s3_c108_n229_c)
    );

    fa fa_s3_c108_n230 (
        .a(stage3_col108[6]),
        .b(stage3_col108[7]),
        .c_in(stage3_col108[8]),
        .s(fa_s3_c108_n230_s),
        .c_out(fa_s3_c108_n230_c)
    );

    fa fa_s3_c109_n231 (
        .a(stage3_col109[0]),
        .b(stage3_col109[1]),
        .c_in(stage3_col109[2]),
        .s(fa_s3_c109_n231_s),
        .c_out(fa_s3_c109_n231_c)
    );

    fa fa_s3_c109_n232 (
        .a(stage3_col109[3]),
        .b(stage3_col109[4]),
        .c_in(stage3_col109[5]),
        .s(fa_s3_c109_n232_s),
        .c_out(fa_s3_c109_n232_c)
    );

    fa fa_s3_c109_n233 (
        .a(stage3_col109[6]),
        .b(stage3_col109[7]),
        .c_in(stage3_col109[8]),
        .s(fa_s3_c109_n233_s),
        .c_out(fa_s3_c109_n233_c)
    );

    fa fa_s3_c110_n234 (
        .a(stage3_col110[0]),
        .b(stage3_col110[1]),
        .c_in(stage3_col110[2]),
        .s(fa_s3_c110_n234_s),
        .c_out(fa_s3_c110_n234_c)
    );

    fa fa_s3_c110_n235 (
        .a(stage3_col110[3]),
        .b(stage3_col110[4]),
        .c_in(stage3_col110[5]),
        .s(fa_s3_c110_n235_s),
        .c_out(fa_s3_c110_n235_c)
    );

    fa fa_s3_c110_n236 (
        .a(stage3_col110[6]),
        .b(stage3_col110[7]),
        .c_in(stage3_col110[8]),
        .s(fa_s3_c110_n236_s),
        .c_out(fa_s3_c110_n236_c)
    );

    fa fa_s3_c111_n237 (
        .a(stage3_col111[0]),
        .b(stage3_col111[1]),
        .c_in(stage3_col111[2]),
        .s(fa_s3_c111_n237_s),
        .c_out(fa_s3_c111_n237_c)
    );

    fa fa_s3_c111_n238 (
        .a(stage3_col111[3]),
        .b(stage3_col111[4]),
        .c_in(stage3_col111[5]),
        .s(fa_s3_c111_n238_s),
        .c_out(fa_s3_c111_n238_c)
    );

    fa fa_s3_c111_n239 (
        .a(stage3_col111[6]),
        .b(stage3_col111[7]),
        .c_in(stage3_col111[8]),
        .s(fa_s3_c111_n239_s),
        .c_out(fa_s3_c111_n239_c)
    );

    fa fa_s3_c112_n240 (
        .a(stage3_col112[0]),
        .b(stage3_col112[1]),
        .c_in(stage3_col112[2]),
        .s(fa_s3_c112_n240_s),
        .c_out(fa_s3_c112_n240_c)
    );

    fa fa_s3_c112_n241 (
        .a(stage3_col112[3]),
        .b(stage3_col112[4]),
        .c_in(stage3_col112[5]),
        .s(fa_s3_c112_n241_s),
        .c_out(fa_s3_c112_n241_c)
    );

    fa fa_s3_c112_n242 (
        .a(stage3_col112[6]),
        .b(stage3_col112[7]),
        .c_in(stage3_col112[8]),
        .s(fa_s3_c112_n242_s),
        .c_out(fa_s3_c112_n242_c)
    );

    fa fa_s3_c113_n243 (
        .a(stage3_col113[0]),
        .b(stage3_col113[1]),
        .c_in(stage3_col113[2]),
        .s(fa_s3_c113_n243_s),
        .c_out(fa_s3_c113_n243_c)
    );

    fa fa_s3_c113_n244 (
        .a(stage3_col113[3]),
        .b(stage3_col113[4]),
        .c_in(stage3_col113[5]),
        .s(fa_s3_c113_n244_s),
        .c_out(fa_s3_c113_n244_c)
    );

    fa fa_s3_c113_n245 (
        .a(stage3_col113[6]),
        .b(stage3_col113[7]),
        .c_in(stage3_col113[8]),
        .s(fa_s3_c113_n245_s),
        .c_out(fa_s3_c113_n245_c)
    );

    fa fa_s3_c114_n246 (
        .a(stage3_col114[0]),
        .b(stage3_col114[1]),
        .c_in(stage3_col114[2]),
        .s(fa_s3_c114_n246_s),
        .c_out(fa_s3_c114_n246_c)
    );

    fa fa_s3_c114_n247 (
        .a(stage3_col114[3]),
        .b(stage3_col114[4]),
        .c_in(stage3_col114[5]),
        .s(fa_s3_c114_n247_s),
        .c_out(fa_s3_c114_n247_c)
    );

    fa fa_s3_c114_n248 (
        .a(stage3_col114[6]),
        .b(stage3_col114[7]),
        .c_in(stage3_col114[8]),
        .s(fa_s3_c114_n248_s),
        .c_out(fa_s3_c114_n248_c)
    );

    fa fa_s3_c115_n249 (
        .a(stage3_col115[0]),
        .b(stage3_col115[1]),
        .c_in(stage3_col115[2]),
        .s(fa_s3_c115_n249_s),
        .c_out(fa_s3_c115_n249_c)
    );

    fa fa_s3_c115_n250 (
        .a(stage3_col115[3]),
        .b(stage3_col115[4]),
        .c_in(stage3_col115[5]),
        .s(fa_s3_c115_n250_s),
        .c_out(fa_s3_c115_n250_c)
    );

    fa fa_s3_c115_n251 (
        .a(stage3_col115[6]),
        .b(stage3_col115[7]),
        .c_in(stage3_col115[8]),
        .s(fa_s3_c115_n251_s),
        .c_out(fa_s3_c115_n251_c)
    );

    fa fa_s3_c116_n252 (
        .a(stage3_col116[0]),
        .b(stage3_col116[1]),
        .c_in(stage3_col116[2]),
        .s(fa_s3_c116_n252_s),
        .c_out(fa_s3_c116_n252_c)
    );

    fa fa_s3_c116_n253 (
        .a(stage3_col116[3]),
        .b(stage3_col116[4]),
        .c_in(stage3_col116[5]),
        .s(fa_s3_c116_n253_s),
        .c_out(fa_s3_c116_n253_c)
    );

    fa fa_s3_c116_n254 (
        .a(stage3_col116[6]),
        .b(stage3_col116[7]),
        .c_in(stage3_col116[8]),
        .s(fa_s3_c116_n254_s),
        .c_out(fa_s3_c116_n254_c)
    );

    fa fa_s3_c117_n255 (
        .a(stage3_col117[0]),
        .b(stage3_col117[1]),
        .c_in(stage3_col117[2]),
        .s(fa_s3_c117_n255_s),
        .c_out(fa_s3_c117_n255_c)
    );

    fa fa_s3_c117_n256 (
        .a(stage3_col117[3]),
        .b(stage3_col117[4]),
        .c_in(stage3_col117[5]),
        .s(fa_s3_c117_n256_s),
        .c_out(fa_s3_c117_n256_c)
    );

    fa fa_s3_c117_n257 (
        .a(stage3_col117[6]),
        .b(stage3_col117[7]),
        .c_in(stage3_col117[8]),
        .s(fa_s3_c117_n257_s),
        .c_out(fa_s3_c117_n257_c)
    );

    fa fa_s3_c118_n258 (
        .a(stage3_col118[0]),
        .b(stage3_col118[1]),
        .c_in(stage3_col118[2]),
        .s(fa_s3_c118_n258_s),
        .c_out(fa_s3_c118_n258_c)
    );

    fa fa_s3_c118_n259 (
        .a(stage3_col118[3]),
        .b(stage3_col118[4]),
        .c_in(stage3_col118[5]),
        .s(fa_s3_c118_n259_s),
        .c_out(fa_s3_c118_n259_c)
    );

    fa fa_s3_c118_n260 (
        .a(stage3_col118[6]),
        .b(stage3_col118[7]),
        .c_in(stage3_col118[8]),
        .s(fa_s3_c118_n260_s),
        .c_out(fa_s3_c118_n260_c)
    );

    fa fa_s3_c119_n261 (
        .a(stage3_col119[0]),
        .b(stage3_col119[1]),
        .c_in(stage3_col119[2]),
        .s(fa_s3_c119_n261_s),
        .c_out(fa_s3_c119_n261_c)
    );

    fa fa_s3_c119_n262 (
        .a(stage3_col119[3]),
        .b(stage3_col119[4]),
        .c_in(stage3_col119[5]),
        .s(fa_s3_c119_n262_s),
        .c_out(fa_s3_c119_n262_c)
    );

    fa fa_s3_c119_n263 (
        .a(stage3_col119[6]),
        .b(stage3_col119[7]),
        .c_in(stage3_col119[8]),
        .s(fa_s3_c119_n263_s),
        .c_out(fa_s3_c119_n263_c)
    );

    fa fa_s3_c120_n264 (
        .a(stage3_col120[0]),
        .b(stage3_col120[1]),
        .c_in(stage3_col120[2]),
        .s(fa_s3_c120_n264_s),
        .c_out(fa_s3_c120_n264_c)
    );

    fa fa_s3_c120_n265 (
        .a(stage3_col120[3]),
        .b(stage3_col120[4]),
        .c_in(stage3_col120[5]),
        .s(fa_s3_c120_n265_s),
        .c_out(fa_s3_c120_n265_c)
    );

    fa fa_s3_c120_n266 (
        .a(stage3_col120[6]),
        .b(stage3_col120[7]),
        .c_in(stage3_col120[8]),
        .s(fa_s3_c120_n266_s),
        .c_out(fa_s3_c120_n266_c)
    );

    fa fa_s3_c121_n267 (
        .a(stage3_col121[0]),
        .b(stage3_col121[1]),
        .c_in(stage3_col121[2]),
        .s(fa_s3_c121_n267_s),
        .c_out(fa_s3_c121_n267_c)
    );

    fa fa_s3_c121_n268 (
        .a(stage3_col121[3]),
        .b(stage3_col121[4]),
        .c_in(stage3_col121[5]),
        .s(fa_s3_c121_n268_s),
        .c_out(fa_s3_c121_n268_c)
    );

    fa fa_s3_c121_n269 (
        .a(stage3_col121[6]),
        .b(stage3_col121[7]),
        .c_in(stage3_col121[8]),
        .s(fa_s3_c121_n269_s),
        .c_out(fa_s3_c121_n269_c)
    );

    fa fa_s3_c122_n270 (
        .a(stage3_col122[0]),
        .b(stage3_col122[1]),
        .c_in(stage3_col122[2]),
        .s(fa_s3_c122_n270_s),
        .c_out(fa_s3_c122_n270_c)
    );

    fa fa_s3_c122_n271 (
        .a(stage3_col122[3]),
        .b(stage3_col122[4]),
        .c_in(stage3_col122[5]),
        .s(fa_s3_c122_n271_s),
        .c_out(fa_s3_c122_n271_c)
    );

    fa fa_s3_c122_n272 (
        .a(stage3_col122[6]),
        .b(stage3_col122[7]),
        .c_in(stage3_col122[8]),
        .s(fa_s3_c122_n272_s),
        .c_out(fa_s3_c122_n272_c)
    );

    fa fa_s3_c123_n273 (
        .a(stage3_col123[0]),
        .b(stage3_col123[1]),
        .c_in(stage3_col123[2]),
        .s(fa_s3_c123_n273_s),
        .c_out(fa_s3_c123_n273_c)
    );

    fa fa_s3_c123_n274 (
        .a(stage3_col123[3]),
        .b(stage3_col123[4]),
        .c_in(stage3_col123[5]),
        .s(fa_s3_c123_n274_s),
        .c_out(fa_s3_c123_n274_c)
    );

    fa fa_s3_c123_n275 (
        .a(stage3_col123[6]),
        .b(stage3_col123[7]),
        .c_in(stage3_col123[8]),
        .s(fa_s3_c123_n275_s),
        .c_out(fa_s3_c123_n275_c)
    );

    fa fa_s3_c124_n276 (
        .a(stage3_col124[0]),
        .b(stage3_col124[1]),
        .c_in(stage3_col124[2]),
        .s(fa_s3_c124_n276_s),
        .c_out(fa_s3_c124_n276_c)
    );

    fa fa_s3_c124_n277 (
        .a(stage3_col124[3]),
        .b(stage3_col124[4]),
        .c_in(stage3_col124[5]),
        .s(fa_s3_c124_n277_s),
        .c_out(fa_s3_c124_n277_c)
    );

    fa fa_s3_c124_n278 (
        .a(stage3_col124[6]),
        .b(stage3_col124[7]),
        .c_in(stage3_col124[8]),
        .s(fa_s3_c124_n278_s),
        .c_out(fa_s3_c124_n278_c)
    );

    fa fa_s3_c125_n279 (
        .a(stage3_col125[0]),
        .b(stage3_col125[1]),
        .c_in(stage3_col125[2]),
        .s(fa_s3_c125_n279_s),
        .c_out(fa_s3_c125_n279_c)
    );

    fa fa_s3_c125_n280 (
        .a(stage3_col125[3]),
        .b(stage3_col125[4]),
        .c_in(stage3_col125[5]),
        .s(fa_s3_c125_n280_s),
        .c_out(fa_s3_c125_n280_c)
    );

    fa fa_s3_c125_n281 (
        .a(stage3_col125[6]),
        .b(stage3_col125[7]),
        .c_in(stage3_col125[8]),
        .s(fa_s3_c125_n281_s),
        .c_out(fa_s3_c125_n281_c)
    );

    fa fa_s3_c126_n282 (
        .a(stage3_col126[0]),
        .b(stage3_col126[1]),
        .c_in(stage3_col126[2]),
        .s(fa_s3_c126_n282_s),
        .c_out(fa_s3_c126_n282_c)
    );

    fa fa_s3_c126_n283 (
        .a(stage3_col126[3]),
        .b(stage3_col126[4]),
        .c_in(stage3_col126[5]),
        .s(fa_s3_c126_n283_s),
        .c_out(fa_s3_c126_n283_c)
    );

    fa fa_s3_c126_n284 (
        .a(stage3_col126[6]),
        .b(stage3_col126[7]),
        .c_in(stage3_col126[8]),
        .s(fa_s3_c126_n284_s),
        .c_out(fa_s3_c126_n284_c)
    );

    ha ha_s3_c3_n0 (
        .a(stage3_col3[0]),
        .b(stage3_col3[1]),
        .s(ha_s3_c3_n0_s),
        .c_out(ha_s3_c3_n0_c)
    );

    // Map to Stage 4 columns
    generate
        if (PIPE) begin : gen_stage4_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage4_col0[0] <= 1'b0;
                    stage4_col1[0] <= 1'b0;
                    stage4_col2[0] <= 1'b0;
                    stage4_col3[0] <= 1'b0;
                    stage4_col4[0] <= 1'b0;
                    stage4_col4[1] <= 1'b0;
                    stage4_col5[0] <= 1'b0;
                    stage4_col6[0] <= 1'b0;
                    stage4_col6[1] <= 1'b0;
                    stage4_col6[2] <= 1'b0;
                    stage4_col7[0] <= 1'b0;
                    stage4_col7[1] <= 1'b0;
                    stage4_col8[0] <= 1'b0;
                    stage4_col8[1] <= 1'b0;
                    stage4_col9[0] <= 1'b0;
                    stage4_col9[1] <= 1'b0;
                    stage4_col10[0] <= 1'b0;
                    stage4_col10[1] <= 1'b0;
                    stage4_col11[0] <= 1'b0;
                    stage4_col11[1] <= 1'b0;
                    stage4_col12[0] <= 1'b0;
                    stage4_col12[1] <= 1'b0;
                    stage4_col13[0] <= 1'b0;
                    stage4_col13[1] <= 1'b0;
                    stage4_col14[0] <= 1'b0;
                    stage4_col14[1] <= 1'b0;
                    stage4_col15[0] <= 1'b0;
                    stage4_col15[1] <= 1'b0;
                    stage4_col16[0] <= 1'b0;
                    stage4_col16[1] <= 1'b0;
                    stage4_col17[0] <= 1'b0;
                    stage4_col17[1] <= 1'b0;
                    stage4_col18[0] <= 1'b0;
                    stage4_col18[1] <= 1'b0;
                    stage4_col19[0] <= 1'b0;
                    stage4_col19[1] <= 1'b0;
                    stage4_col19[2] <= 1'b0;
                    stage4_col19[3] <= 1'b0;
                    stage4_col20[0] <= 1'b0;
                    stage4_col20[1] <= 1'b0;
                    stage4_col20[2] <= 1'b0;
                    stage4_col21[0] <= 1'b0;
                    stage4_col21[1] <= 1'b0;
                    stage4_col21[2] <= 1'b0;
                    stage4_col22[0] <= 1'b0;
                    stage4_col22[1] <= 1'b0;
                    stage4_col22[2] <= 1'b0;
                    stage4_col23[0] <= 1'b0;
                    stage4_col23[1] <= 1'b0;
                    stage4_col23[2] <= 1'b0;
                    stage4_col24[0] <= 1'b0;
                    stage4_col24[1] <= 1'b0;
                    stage4_col24[2] <= 1'b0;
                    stage4_col25[0] <= 1'b0;
                    stage4_col25[1] <= 1'b0;
                    stage4_col25[2] <= 1'b0;
                    stage4_col26[0] <= 1'b0;
                    stage4_col26[1] <= 1'b0;
                    stage4_col26[2] <= 1'b0;
                    stage4_col27[0] <= 1'b0;
                    stage4_col27[1] <= 1'b0;
                    stage4_col27[2] <= 1'b0;
                    stage4_col28[0] <= 1'b0;
                    stage4_col28[1] <= 1'b0;
                    stage4_col28[2] <= 1'b0;
                    stage4_col28[3] <= 1'b0;
                    stage4_col28[4] <= 1'b0;
                    stage4_col29[0] <= 1'b0;
                    stage4_col29[1] <= 1'b0;
                    stage4_col29[2] <= 1'b0;
                    stage4_col29[3] <= 1'b0;
                    stage4_col30[0] <= 1'b0;
                    stage4_col30[1] <= 1'b0;
                    stage4_col30[2] <= 1'b0;
                    stage4_col30[3] <= 1'b0;
                    stage4_col31[0] <= 1'b0;
                    stage4_col31[1] <= 1'b0;
                    stage4_col31[2] <= 1'b0;
                    stage4_col31[3] <= 1'b0;
                    stage4_col32[0] <= 1'b0;
                    stage4_col32[1] <= 1'b0;
                    stage4_col32[2] <= 1'b0;
                    stage4_col32[3] <= 1'b0;
                    stage4_col33[0] <= 1'b0;
                    stage4_col33[1] <= 1'b0;
                    stage4_col33[2] <= 1'b0;
                    stage4_col33[3] <= 1'b0;
                    stage4_col34[0] <= 1'b0;
                    stage4_col34[1] <= 1'b0;
                    stage4_col34[2] <= 1'b0;
                    stage4_col34[3] <= 1'b0;
                    stage4_col35[0] <= 1'b0;
                    stage4_col35[1] <= 1'b0;
                    stage4_col35[2] <= 1'b0;
                    stage4_col35[3] <= 1'b0;
                    stage4_col36[0] <= 1'b0;
                    stage4_col36[1] <= 1'b0;
                    stage4_col36[2] <= 1'b0;
                    stage4_col36[3] <= 1'b0;
                    stage4_col37[0] <= 1'b0;
                    stage4_col37[1] <= 1'b0;
                    stage4_col37[2] <= 1'b0;
                    stage4_col37[3] <= 1'b0;
                    stage4_col38[0] <= 1'b0;
                    stage4_col38[1] <= 1'b0;
                    stage4_col38[2] <= 1'b0;
                    stage4_col38[3] <= 1'b0;
                    stage4_col39[0] <= 1'b0;
                    stage4_col39[1] <= 1'b0;
                    stage4_col39[2] <= 1'b0;
                    stage4_col39[3] <= 1'b0;
                    stage4_col40[0] <= 1'b0;
                    stage4_col40[1] <= 1'b0;
                    stage4_col40[2] <= 1'b0;
                    stage4_col40[3] <= 1'b0;
                    stage4_col40[4] <= 1'b0;
                    stage4_col40[5] <= 1'b0;
                    stage4_col41[0] <= 1'b0;
                    stage4_col41[1] <= 1'b0;
                    stage4_col41[2] <= 1'b0;
                    stage4_col41[3] <= 1'b0;
                    stage4_col41[4] <= 1'b0;
                    stage4_col42[0] <= 1'b0;
                    stage4_col42[1] <= 1'b0;
                    stage4_col42[2] <= 1'b0;
                    stage4_col42[3] <= 1'b0;
                    stage4_col42[4] <= 1'b0;
                    stage4_col43[0] <= 1'b0;
                    stage4_col43[1] <= 1'b0;
                    stage4_col43[2] <= 1'b0;
                    stage4_col43[3] <= 1'b0;
                    stage4_col43[4] <= 1'b0;
                    stage4_col44[0] <= 1'b0;
                    stage4_col44[1] <= 1'b0;
                    stage4_col44[2] <= 1'b0;
                    stage4_col44[3] <= 1'b0;
                    stage4_col44[4] <= 1'b0;
                    stage4_col45[0] <= 1'b0;
                    stage4_col45[1] <= 1'b0;
                    stage4_col45[2] <= 1'b0;
                    stage4_col45[3] <= 1'b0;
                    stage4_col45[4] <= 1'b0;
                    stage4_col46[0] <= 1'b0;
                    stage4_col46[1] <= 1'b0;
                    stage4_col46[2] <= 1'b0;
                    stage4_col46[3] <= 1'b0;
                    stage4_col46[4] <= 1'b0;
                    stage4_col47[0] <= 1'b0;
                    stage4_col47[1] <= 1'b0;
                    stage4_col47[2] <= 1'b0;
                    stage4_col47[3] <= 1'b0;
                    stage4_col47[4] <= 1'b0;
                    stage4_col47[5] <= 1'b0;
                    stage4_col47[6] <= 1'b0;
                    stage4_col48[0] <= 1'b0;
                    stage4_col48[1] <= 1'b0;
                    stage4_col48[2] <= 1'b0;
                    stage4_col48[3] <= 1'b0;
                    stage4_col48[4] <= 1'b0;
                    stage4_col48[5] <= 1'b0;
                    stage4_col49[0] <= 1'b0;
                    stage4_col49[1] <= 1'b0;
                    stage4_col49[2] <= 1'b0;
                    stage4_col49[3] <= 1'b0;
                    stage4_col49[4] <= 1'b0;
                    stage4_col49[5] <= 1'b0;
                    stage4_col50[0] <= 1'b0;
                    stage4_col50[1] <= 1'b0;
                    stage4_col50[2] <= 1'b0;
                    stage4_col50[3] <= 1'b0;
                    stage4_col50[4] <= 1'b0;
                    stage4_col50[5] <= 1'b0;
                    stage4_col51[0] <= 1'b0;
                    stage4_col51[1] <= 1'b0;
                    stage4_col51[2] <= 1'b0;
                    stage4_col51[3] <= 1'b0;
                    stage4_col51[4] <= 1'b0;
                    stage4_col51[5] <= 1'b0;
                    stage4_col52[0] <= 1'b0;
                    stage4_col52[1] <= 1'b0;
                    stage4_col52[2] <= 1'b0;
                    stage4_col52[3] <= 1'b0;
                    stage4_col52[4] <= 1'b0;
                    stage4_col52[5] <= 1'b0;
                    stage4_col53[0] <= 1'b0;
                    stage4_col53[1] <= 1'b0;
                    stage4_col53[2] <= 1'b0;
                    stage4_col53[3] <= 1'b0;
                    stage4_col53[4] <= 1'b0;
                    stage4_col53[5] <= 1'b0;
                    stage4_col54[0] <= 1'b0;
                    stage4_col54[1] <= 1'b0;
                    stage4_col54[2] <= 1'b0;
                    stage4_col54[3] <= 1'b0;
                    stage4_col54[4] <= 1'b0;
                    stage4_col54[5] <= 1'b0;
                    stage4_col55[0] <= 1'b0;
                    stage4_col55[1] <= 1'b0;
                    stage4_col55[2] <= 1'b0;
                    stage4_col55[3] <= 1'b0;
                    stage4_col55[4] <= 1'b0;
                    stage4_col55[5] <= 1'b0;
                    stage4_col56[0] <= 1'b0;
                    stage4_col56[1] <= 1'b0;
                    stage4_col56[2] <= 1'b0;
                    stage4_col56[3] <= 1'b0;
                    stage4_col56[4] <= 1'b0;
                    stage4_col56[5] <= 1'b0;
                    stage4_col57[0] <= 1'b0;
                    stage4_col57[1] <= 1'b0;
                    stage4_col57[2] <= 1'b0;
                    stage4_col57[3] <= 1'b0;
                    stage4_col57[4] <= 1'b0;
                    stage4_col57[5] <= 1'b0;
                    stage4_col58[0] <= 1'b0;
                    stage4_col58[1] <= 1'b0;
                    stage4_col58[2] <= 1'b0;
                    stage4_col58[3] <= 1'b0;
                    stage4_col58[4] <= 1'b0;
                    stage4_col58[5] <= 1'b0;
                    stage4_col59[0] <= 1'b0;
                    stage4_col59[1] <= 1'b0;
                    stage4_col59[2] <= 1'b0;
                    stage4_col59[3] <= 1'b0;
                    stage4_col59[4] <= 1'b0;
                    stage4_col59[5] <= 1'b0;
                    stage4_col59[6] <= 1'b0;
                    stage4_col59[7] <= 1'b0;
                    stage4_col60[0] <= 1'b0;
                    stage4_col60[1] <= 1'b0;
                    stage4_col60[2] <= 1'b0;
                    stage4_col60[3] <= 1'b0;
                    stage4_col60[4] <= 1'b0;
                    stage4_col60[5] <= 1'b0;
                    stage4_col60[6] <= 1'b0;
                    stage4_col61[0] <= 1'b0;
                    stage4_col61[1] <= 1'b0;
                    stage4_col61[2] <= 1'b0;
                    stage4_col61[3] <= 1'b0;
                    stage4_col61[4] <= 1'b0;
                    stage4_col61[5] <= 1'b0;
                    stage4_col61[6] <= 1'b0;
                    stage4_col62[0] <= 1'b0;
                    stage4_col62[1] <= 1'b0;
                    stage4_col62[2] <= 1'b0;
                    stage4_col62[3] <= 1'b0;
                    stage4_col62[4] <= 1'b0;
                    stage4_col62[5] <= 1'b0;
                    stage4_col62[6] <= 1'b0;
                    stage4_col63[0] <= 1'b0;
                    stage4_col63[1] <= 1'b0;
                    stage4_col63[2] <= 1'b0;
                    stage4_col63[3] <= 1'b0;
                    stage4_col63[4] <= 1'b0;
                    stage4_col63[5] <= 1'b0;
                    stage4_col63[6] <= 1'b0;
                    stage4_col64[0] <= 1'b0;
                    stage4_col64[1] <= 1'b0;
                    stage4_col64[2] <= 1'b0;
                    stage4_col64[3] <= 1'b0;
                    stage4_col64[4] <= 1'b0;
                    stage4_col64[5] <= 1'b0;
                    stage4_col64[6] <= 1'b0;
                    stage4_col64[7] <= 1'b0;
                    stage4_col65[0] <= 1'b0;
                    stage4_col65[1] <= 1'b0;
                    stage4_col65[2] <= 1'b0;
                    stage4_col65[3] <= 1'b0;
                    stage4_col65[4] <= 1'b0;
                    stage4_col65[5] <= 1'b0;
                    stage4_col65[6] <= 1'b0;
                    stage4_col66[0] <= 1'b0;
                    stage4_col66[1] <= 1'b0;
                    stage4_col66[2] <= 1'b0;
                    stage4_col66[3] <= 1'b0;
                    stage4_col66[4] <= 1'b0;
                    stage4_col66[5] <= 1'b0;
                    stage4_col66[6] <= 1'b0;
                    stage4_col66[7] <= 1'b0;
                    stage4_col67[0] <= 1'b0;
                    stage4_col67[1] <= 1'b0;
                    stage4_col67[2] <= 1'b0;
                    stage4_col67[3] <= 1'b0;
                    stage4_col67[4] <= 1'b0;
                    stage4_col67[5] <= 1'b0;
                    stage4_col67[6] <= 1'b0;
                    stage4_col68[0] <= 1'b0;
                    stage4_col68[1] <= 1'b0;
                    stage4_col68[2] <= 1'b0;
                    stage4_col68[3] <= 1'b0;
                    stage4_col68[4] <= 1'b0;
                    stage4_col68[5] <= 1'b0;
                    stage4_col68[6] <= 1'b0;
                    stage4_col68[7] <= 1'b0;
                    stage4_col69[0] <= 1'b0;
                    stage4_col69[1] <= 1'b0;
                    stage4_col69[2] <= 1'b0;
                    stage4_col69[3] <= 1'b0;
                    stage4_col69[4] <= 1'b0;
                    stage4_col69[5] <= 1'b0;
                    stage4_col69[6] <= 1'b0;
                    stage4_col70[0] <= 1'b0;
                    stage4_col70[1] <= 1'b0;
                    stage4_col70[2] <= 1'b0;
                    stage4_col70[3] <= 1'b0;
                    stage4_col70[4] <= 1'b0;
                    stage4_col70[5] <= 1'b0;
                    stage4_col70[6] <= 1'b0;
                    stage4_col70[7] <= 1'b0;
                    stage4_col71[0] <= 1'b0;
                    stage4_col71[1] <= 1'b0;
                    stage4_col71[2] <= 1'b0;
                    stage4_col71[3] <= 1'b0;
                    stage4_col71[4] <= 1'b0;
                    stage4_col71[5] <= 1'b0;
                    stage4_col71[6] <= 1'b0;
                    stage4_col72[0] <= 1'b0;
                    stage4_col72[1] <= 1'b0;
                    stage4_col72[2] <= 1'b0;
                    stage4_col72[3] <= 1'b0;
                    stage4_col72[4] <= 1'b0;
                    stage4_col72[5] <= 1'b0;
                    stage4_col72[6] <= 1'b0;
                    stage4_col72[7] <= 1'b0;
                    stage4_col73[0] <= 1'b0;
                    stage4_col73[1] <= 1'b0;
                    stage4_col73[2] <= 1'b0;
                    stage4_col73[3] <= 1'b0;
                    stage4_col73[4] <= 1'b0;
                    stage4_col73[5] <= 1'b0;
                    stage4_col73[6] <= 1'b0;
                    stage4_col74[0] <= 1'b0;
                    stage4_col74[1] <= 1'b0;
                    stage4_col74[2] <= 1'b0;
                    stage4_col74[3] <= 1'b0;
                    stage4_col74[4] <= 1'b0;
                    stage4_col74[5] <= 1'b0;
                    stage4_col74[6] <= 1'b0;
                    stage4_col74[7] <= 1'b0;
                    stage4_col75[0] <= 1'b0;
                    stage4_col75[1] <= 1'b0;
                    stage4_col75[2] <= 1'b0;
                    stage4_col75[3] <= 1'b0;
                    stage4_col75[4] <= 1'b0;
                    stage4_col75[5] <= 1'b0;
                    stage4_col75[6] <= 1'b0;
                    stage4_col76[0] <= 1'b0;
                    stage4_col76[1] <= 1'b0;
                    stage4_col76[2] <= 1'b0;
                    stage4_col76[3] <= 1'b0;
                    stage4_col76[4] <= 1'b0;
                    stage4_col76[5] <= 1'b0;
                    stage4_col76[6] <= 1'b0;
                    stage4_col76[7] <= 1'b0;
                    stage4_col77[0] <= 1'b0;
                    stage4_col77[1] <= 1'b0;
                    stage4_col77[2] <= 1'b0;
                    stage4_col77[3] <= 1'b0;
                    stage4_col77[4] <= 1'b0;
                    stage4_col77[5] <= 1'b0;
                    stage4_col77[6] <= 1'b0;
                    stage4_col78[0] <= 1'b0;
                    stage4_col78[1] <= 1'b0;
                    stage4_col78[2] <= 1'b0;
                    stage4_col78[3] <= 1'b0;
                    stage4_col78[4] <= 1'b0;
                    stage4_col78[5] <= 1'b0;
                    stage4_col78[6] <= 1'b0;
                    stage4_col78[7] <= 1'b0;
                    stage4_col79[0] <= 1'b0;
                    stage4_col79[1] <= 1'b0;
                    stage4_col79[2] <= 1'b0;
                    stage4_col79[3] <= 1'b0;
                    stage4_col79[4] <= 1'b0;
                    stage4_col79[5] <= 1'b0;
                    stage4_col79[6] <= 1'b0;
                    stage4_col80[0] <= 1'b0;
                    stage4_col80[1] <= 1'b0;
                    stage4_col80[2] <= 1'b0;
                    stage4_col80[3] <= 1'b0;
                    stage4_col80[4] <= 1'b0;
                    stage4_col80[5] <= 1'b0;
                    stage4_col80[6] <= 1'b0;
                    stage4_col80[7] <= 1'b0;
                    stage4_col81[0] <= 1'b0;
                    stage4_col81[1] <= 1'b0;
                    stage4_col81[2] <= 1'b0;
                    stage4_col81[3] <= 1'b0;
                    stage4_col81[4] <= 1'b0;
                    stage4_col81[5] <= 1'b0;
                    stage4_col81[6] <= 1'b0;
                    stage4_col82[0] <= 1'b0;
                    stage4_col82[1] <= 1'b0;
                    stage4_col82[2] <= 1'b0;
                    stage4_col82[3] <= 1'b0;
                    stage4_col82[4] <= 1'b0;
                    stage4_col82[5] <= 1'b0;
                    stage4_col82[6] <= 1'b0;
                    stage4_col82[7] <= 1'b0;
                    stage4_col83[0] <= 1'b0;
                    stage4_col83[1] <= 1'b0;
                    stage4_col83[2] <= 1'b0;
                    stage4_col83[3] <= 1'b0;
                    stage4_col83[4] <= 1'b0;
                    stage4_col83[5] <= 1'b0;
                    stage4_col83[6] <= 1'b0;
                    stage4_col84[0] <= 1'b0;
                    stage4_col84[1] <= 1'b0;
                    stage4_col84[2] <= 1'b0;
                    stage4_col84[3] <= 1'b0;
                    stage4_col84[4] <= 1'b0;
                    stage4_col84[5] <= 1'b0;
                    stage4_col84[6] <= 1'b0;
                    stage4_col84[7] <= 1'b0;
                    stage4_col85[0] <= 1'b0;
                    stage4_col85[1] <= 1'b0;
                    stage4_col85[2] <= 1'b0;
                    stage4_col85[3] <= 1'b0;
                    stage4_col85[4] <= 1'b0;
                    stage4_col85[5] <= 1'b0;
                    stage4_col85[6] <= 1'b0;
                    stage4_col86[0] <= 1'b0;
                    stage4_col86[1] <= 1'b0;
                    stage4_col86[2] <= 1'b0;
                    stage4_col86[3] <= 1'b0;
                    stage4_col86[4] <= 1'b0;
                    stage4_col86[5] <= 1'b0;
                    stage4_col86[6] <= 1'b0;
                    stage4_col86[7] <= 1'b0;
                    stage4_col87[0] <= 1'b0;
                    stage4_col87[1] <= 1'b0;
                    stage4_col87[2] <= 1'b0;
                    stage4_col87[3] <= 1'b0;
                    stage4_col87[4] <= 1'b0;
                    stage4_col87[5] <= 1'b0;
                    stage4_col87[6] <= 1'b0;
                    stage4_col88[0] <= 1'b0;
                    stage4_col88[1] <= 1'b0;
                    stage4_col88[2] <= 1'b0;
                    stage4_col88[3] <= 1'b0;
                    stage4_col88[4] <= 1'b0;
                    stage4_col88[5] <= 1'b0;
                    stage4_col88[6] <= 1'b0;
                    stage4_col88[7] <= 1'b0;
                    stage4_col89[0] <= 1'b0;
                    stage4_col89[1] <= 1'b0;
                    stage4_col89[2] <= 1'b0;
                    stage4_col89[3] <= 1'b0;
                    stage4_col89[4] <= 1'b0;
                    stage4_col89[5] <= 1'b0;
                    stage4_col89[6] <= 1'b0;
                    stage4_col90[0] <= 1'b0;
                    stage4_col90[1] <= 1'b0;
                    stage4_col90[2] <= 1'b0;
                    stage4_col90[3] <= 1'b0;
                    stage4_col90[4] <= 1'b0;
                    stage4_col90[5] <= 1'b0;
                    stage4_col90[6] <= 1'b0;
                    stage4_col90[7] <= 1'b0;
                    stage4_col91[0] <= 1'b0;
                    stage4_col91[1] <= 1'b0;
                    stage4_col91[2] <= 1'b0;
                    stage4_col91[3] <= 1'b0;
                    stage4_col91[4] <= 1'b0;
                    stage4_col91[5] <= 1'b0;
                    stage4_col91[6] <= 1'b0;
                    stage4_col92[0] <= 1'b0;
                    stage4_col92[1] <= 1'b0;
                    stage4_col92[2] <= 1'b0;
                    stage4_col92[3] <= 1'b0;
                    stage4_col92[4] <= 1'b0;
                    stage4_col92[5] <= 1'b0;
                    stage4_col92[6] <= 1'b0;
                    stage4_col92[7] <= 1'b0;
                    stage4_col93[0] <= 1'b0;
                    stage4_col93[1] <= 1'b0;
                    stage4_col93[2] <= 1'b0;
                    stage4_col93[3] <= 1'b0;
                    stage4_col93[4] <= 1'b0;
                    stage4_col93[5] <= 1'b0;
                    stage4_col93[6] <= 1'b0;
                    stage4_col94[0] <= 1'b0;
                    stage4_col94[1] <= 1'b0;
                    stage4_col94[2] <= 1'b0;
                    stage4_col94[3] <= 1'b0;
                    stage4_col94[4] <= 1'b0;
                    stage4_col94[5] <= 1'b0;
                    stage4_col94[6] <= 1'b0;
                    stage4_col94[7] <= 1'b0;
                    stage4_col95[0] <= 1'b0;
                    stage4_col95[1] <= 1'b0;
                    stage4_col95[2] <= 1'b0;
                    stage4_col95[3] <= 1'b0;
                    stage4_col95[4] <= 1'b0;
                    stage4_col95[5] <= 1'b0;
                    stage4_col95[6] <= 1'b0;
                    stage4_col96[0] <= 1'b0;
                    stage4_col96[1] <= 1'b0;
                    stage4_col96[2] <= 1'b0;
                    stage4_col96[3] <= 1'b0;
                    stage4_col96[4] <= 1'b0;
                    stage4_col96[5] <= 1'b0;
                    stage4_col96[6] <= 1'b0;
                    stage4_col96[7] <= 1'b0;
                    stage4_col97[0] <= 1'b0;
                    stage4_col97[1] <= 1'b0;
                    stage4_col97[2] <= 1'b0;
                    stage4_col97[3] <= 1'b0;
                    stage4_col97[4] <= 1'b0;
                    stage4_col97[5] <= 1'b0;
                    stage4_col97[6] <= 1'b0;
                    stage4_col98[0] <= 1'b0;
                    stage4_col98[1] <= 1'b0;
                    stage4_col98[2] <= 1'b0;
                    stage4_col98[3] <= 1'b0;
                    stage4_col98[4] <= 1'b0;
                    stage4_col98[5] <= 1'b0;
                    stage4_col98[6] <= 1'b0;
                    stage4_col98[7] <= 1'b0;
                    stage4_col99[0] <= 1'b0;
                    stage4_col99[1] <= 1'b0;
                    stage4_col99[2] <= 1'b0;
                    stage4_col99[3] <= 1'b0;
                    stage4_col99[4] <= 1'b0;
                    stage4_col99[5] <= 1'b0;
                    stage4_col99[6] <= 1'b0;
                    stage4_col100[0] <= 1'b0;
                    stage4_col100[1] <= 1'b0;
                    stage4_col100[2] <= 1'b0;
                    stage4_col100[3] <= 1'b0;
                    stage4_col100[4] <= 1'b0;
                    stage4_col100[5] <= 1'b0;
                    stage4_col100[6] <= 1'b0;
                    stage4_col100[7] <= 1'b0;
                    stage4_col101[0] <= 1'b0;
                    stage4_col101[1] <= 1'b0;
                    stage4_col101[2] <= 1'b0;
                    stage4_col101[3] <= 1'b0;
                    stage4_col101[4] <= 1'b0;
                    stage4_col101[5] <= 1'b0;
                    stage4_col101[6] <= 1'b0;
                    stage4_col102[0] <= 1'b0;
                    stage4_col102[1] <= 1'b0;
                    stage4_col102[2] <= 1'b0;
                    stage4_col102[3] <= 1'b0;
                    stage4_col102[4] <= 1'b0;
                    stage4_col102[5] <= 1'b0;
                    stage4_col102[6] <= 1'b0;
                    stage4_col102[7] <= 1'b0;
                    stage4_col103[0] <= 1'b0;
                    stage4_col103[1] <= 1'b0;
                    stage4_col103[2] <= 1'b0;
                    stage4_col103[3] <= 1'b0;
                    stage4_col103[4] <= 1'b0;
                    stage4_col103[5] <= 1'b0;
                    stage4_col103[6] <= 1'b0;
                    stage4_col104[0] <= 1'b0;
                    stage4_col104[1] <= 1'b0;
                    stage4_col104[2] <= 1'b0;
                    stage4_col104[3] <= 1'b0;
                    stage4_col104[4] <= 1'b0;
                    stage4_col104[5] <= 1'b0;
                    stage4_col104[6] <= 1'b0;
                    stage4_col104[7] <= 1'b0;
                    stage4_col105[0] <= 1'b0;
                    stage4_col105[1] <= 1'b0;
                    stage4_col105[2] <= 1'b0;
                    stage4_col105[3] <= 1'b0;
                    stage4_col105[4] <= 1'b0;
                    stage4_col105[5] <= 1'b0;
                    stage4_col105[6] <= 1'b0;
                    stage4_col106[0] <= 1'b0;
                    stage4_col106[1] <= 1'b0;
                    stage4_col106[2] <= 1'b0;
                    stage4_col106[3] <= 1'b0;
                    stage4_col106[4] <= 1'b0;
                    stage4_col106[5] <= 1'b0;
                    stage4_col106[6] <= 1'b0;
                    stage4_col106[7] <= 1'b0;
                    stage4_col107[0] <= 1'b0;
                    stage4_col107[1] <= 1'b0;
                    stage4_col107[2] <= 1'b0;
                    stage4_col107[3] <= 1'b0;
                    stage4_col107[4] <= 1'b0;
                    stage4_col107[5] <= 1'b0;
                    stage4_col107[6] <= 1'b0;
                    stage4_col108[0] <= 1'b0;
                    stage4_col108[1] <= 1'b0;
                    stage4_col108[2] <= 1'b0;
                    stage4_col108[3] <= 1'b0;
                    stage4_col108[4] <= 1'b0;
                    stage4_col108[5] <= 1'b0;
                    stage4_col108[6] <= 1'b0;
                    stage4_col108[7] <= 1'b0;
                    stage4_col109[0] <= 1'b0;
                    stage4_col109[1] <= 1'b0;
                    stage4_col109[2] <= 1'b0;
                    stage4_col109[3] <= 1'b0;
                    stage4_col109[4] <= 1'b0;
                    stage4_col109[5] <= 1'b0;
                    stage4_col109[6] <= 1'b0;
                    stage4_col110[0] <= 1'b0;
                    stage4_col110[1] <= 1'b0;
                    stage4_col110[2] <= 1'b0;
                    stage4_col110[3] <= 1'b0;
                    stage4_col110[4] <= 1'b0;
                    stage4_col110[5] <= 1'b0;
                    stage4_col110[6] <= 1'b0;
                    stage4_col110[7] <= 1'b0;
                    stage4_col111[0] <= 1'b0;
                    stage4_col111[1] <= 1'b0;
                    stage4_col111[2] <= 1'b0;
                    stage4_col111[3] <= 1'b0;
                    stage4_col111[4] <= 1'b0;
                    stage4_col111[5] <= 1'b0;
                    stage4_col111[6] <= 1'b0;
                    stage4_col112[0] <= 1'b0;
                    stage4_col112[1] <= 1'b0;
                    stage4_col112[2] <= 1'b0;
                    stage4_col112[3] <= 1'b0;
                    stage4_col112[4] <= 1'b0;
                    stage4_col112[5] <= 1'b0;
                    stage4_col112[6] <= 1'b0;
                    stage4_col112[7] <= 1'b0;
                    stage4_col113[0] <= 1'b0;
                    stage4_col113[1] <= 1'b0;
                    stage4_col113[2] <= 1'b0;
                    stage4_col113[3] <= 1'b0;
                    stage4_col113[4] <= 1'b0;
                    stage4_col113[5] <= 1'b0;
                    stage4_col113[6] <= 1'b0;
                    stage4_col114[0] <= 1'b0;
                    stage4_col114[1] <= 1'b0;
                    stage4_col114[2] <= 1'b0;
                    stage4_col114[3] <= 1'b0;
                    stage4_col114[4] <= 1'b0;
                    stage4_col114[5] <= 1'b0;
                    stage4_col114[6] <= 1'b0;
                    stage4_col114[7] <= 1'b0;
                    stage4_col115[0] <= 1'b0;
                    stage4_col115[1] <= 1'b0;
                    stage4_col115[2] <= 1'b0;
                    stage4_col115[3] <= 1'b0;
                    stage4_col115[4] <= 1'b0;
                    stage4_col115[5] <= 1'b0;
                    stage4_col115[6] <= 1'b0;
                    stage4_col116[0] <= 1'b0;
                    stage4_col116[1] <= 1'b0;
                    stage4_col116[2] <= 1'b0;
                    stage4_col116[3] <= 1'b0;
                    stage4_col116[4] <= 1'b0;
                    stage4_col116[5] <= 1'b0;
                    stage4_col116[6] <= 1'b0;
                    stage4_col116[7] <= 1'b0;
                    stage4_col117[0] <= 1'b0;
                    stage4_col117[1] <= 1'b0;
                    stage4_col117[2] <= 1'b0;
                    stage4_col117[3] <= 1'b0;
                    stage4_col117[4] <= 1'b0;
                    stage4_col117[5] <= 1'b0;
                    stage4_col117[6] <= 1'b0;
                    stage4_col118[0] <= 1'b0;
                    stage4_col118[1] <= 1'b0;
                    stage4_col118[2] <= 1'b0;
                    stage4_col118[3] <= 1'b0;
                    stage4_col118[4] <= 1'b0;
                    stage4_col118[5] <= 1'b0;
                    stage4_col118[6] <= 1'b0;
                    stage4_col118[7] <= 1'b0;
                    stage4_col119[0] <= 1'b0;
                    stage4_col119[1] <= 1'b0;
                    stage4_col119[2] <= 1'b0;
                    stage4_col119[3] <= 1'b0;
                    stage4_col119[4] <= 1'b0;
                    stage4_col119[5] <= 1'b0;
                    stage4_col119[6] <= 1'b0;
                    stage4_col120[0] <= 1'b0;
                    stage4_col120[1] <= 1'b0;
                    stage4_col120[2] <= 1'b0;
                    stage4_col120[3] <= 1'b0;
                    stage4_col120[4] <= 1'b0;
                    stage4_col120[5] <= 1'b0;
                    stage4_col120[6] <= 1'b0;
                    stage4_col120[7] <= 1'b0;
                    stage4_col121[0] <= 1'b0;
                    stage4_col121[1] <= 1'b0;
                    stage4_col121[2] <= 1'b0;
                    stage4_col121[3] <= 1'b0;
                    stage4_col121[4] <= 1'b0;
                    stage4_col121[5] <= 1'b0;
                    stage4_col121[6] <= 1'b0;
                    stage4_col122[0] <= 1'b0;
                    stage4_col122[1] <= 1'b0;
                    stage4_col122[2] <= 1'b0;
                    stage4_col122[3] <= 1'b0;
                    stage4_col122[4] <= 1'b0;
                    stage4_col122[5] <= 1'b0;
                    stage4_col122[6] <= 1'b0;
                    stage4_col122[7] <= 1'b0;
                    stage4_col123[0] <= 1'b0;
                    stage4_col123[1] <= 1'b0;
                    stage4_col123[2] <= 1'b0;
                    stage4_col123[3] <= 1'b0;
                    stage4_col123[4] <= 1'b0;
                    stage4_col123[5] <= 1'b0;
                    stage4_col123[6] <= 1'b0;
                    stage4_col124[0] <= 1'b0;
                    stage4_col124[1] <= 1'b0;
                    stage4_col124[2] <= 1'b0;
                    stage4_col124[3] <= 1'b0;
                    stage4_col124[4] <= 1'b0;
                    stage4_col124[5] <= 1'b0;
                    stage4_col124[6] <= 1'b0;
                    stage4_col124[7] <= 1'b0;
                    stage4_col125[0] <= 1'b0;
                    stage4_col125[1] <= 1'b0;
                    stage4_col125[2] <= 1'b0;
                    stage4_col125[3] <= 1'b0;
                    stage4_col125[4] <= 1'b0;
                    stage4_col125[5] <= 1'b0;
                    stage4_col125[6] <= 1'b0;
                    stage4_col126[0] <= 1'b0;
                    stage4_col126[1] <= 1'b0;
                    stage4_col126[2] <= 1'b0;
                    stage4_col126[3] <= 1'b0;
                    stage4_col126[4] <= 1'b0;
                    stage4_col126[5] <= 1'b0;
                    stage4_col126[6] <= 1'b0;
                    stage4_col126[7] <= 1'b0;
                    stage4_col127[0] <= 1'b0;
                    stage4_col127[1] <= 1'b0;
                    stage4_col127[2] <= 1'b0;
                    stage4_col127[3] <= 1'b0;
                    stage4_col127[4] <= 1'b0;
                    stage4_col127[5] <= 1'b0;
                    stage4_col127[6] <= 1'b0;
                    stage4_col127[7] <= 1'b0;
                    stage4_col127[8] <= 1'b0;
                    stage4_col127[9] <= 1'b0;
                    stage4_col127[10] <= 1'b0;
                    stage4_col127[11] <= 1'b0;
                    stage4_col127[12] <= 1'b0;
                    stage4_col127[13] <= 1'b0;
                    stage4_col127[14] <= 1'b0;
                    stage4_col127[15] <= 1'b0;
                    stage4_col127[16] <= 1'b0;
                    stage4_col127[17] <= 1'b0;
                    stage4_col127[18] <= 1'b0;
                    stage4_col127[19] <= 1'b0;
                    stage4_col127[20] <= 1'b0;
                    stage4_col127[21] <= 1'b0;
                    stage4_col127[22] <= 1'b0;
                    stage4_col127[23] <= 1'b0;
                    stage4_col127[24] <= 1'b0;
                    stage4_col127[25] <= 1'b0;
                    stage4_col127[26] <= 1'b0;
                    stage4_col127[27] <= 1'b0;
                    stage4_col127[28] <= 1'b0;
                    stage4_col127[29] <= 1'b0;
                    stage4_col127[30] <= 1'b0;
                    stage4_col127[31] <= 1'b0;
                    stage4_col127[32] <= 1'b0;
                    stage4_col127[33] <= 1'b0;
                    stage4_col127[34] <= 1'b0;
                    stage4_col127[35] <= 1'b0;
                    stage4_col127[36] <= 1'b0;
                    stage4_col127[37] <= 1'b0;
                    stage4_col127[38] <= 1'b0;
                    stage4_col127[39] <= 1'b0;
                    stage4_col127[40] <= 1'b0;
                    stage4_col127[41] <= 1'b0;
                    stage4_col127[42] <= 1'b0;
                    stage4_col127[43] <= 1'b0;
                    stage4_col127[44] <= 1'b0;
                    stage4_col127[45] <= 1'b0;
                    stage4_col127[46] <= 1'b0;
                    stage4_col127[47] <= 1'b0;
                    stage4_col127[48] <= 1'b0;
                    stage4_col127[49] <= 1'b0;
                    stage4_col127[50] <= 1'b0;
                    stage4_col127[51] <= 1'b0;
                    stage4_col127[52] <= 1'b0;
                    stage4_col127[53] <= 1'b0;
                    stage4_col127[54] <= 1'b0;
                    stage4_col127[55] <= 1'b0;
                    stage4_col127[56] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage4_col0[0] <= stage3_col0[0];
                    stage4_col1[0] <= stage3_col1[0];
                    stage4_col2[0] <= stage3_col2[0];
                    stage4_col3[0] <= ha_s3_c3_n0_s;
                    stage4_col4[0] <= ha_s3_c3_n0_c;
                    stage4_col4[1] <= stage3_col4[0];
                    stage4_col5[0] <= fa_s3_c5_n0_s;
                    stage4_col6[0] <= fa_s3_c5_n0_c;
                    stage4_col6[1] <= stage3_col6[0];
                    stage4_col6[2] <= stage3_col6[1];
                    stage4_col7[0] <= stage3_col7[0];
                    stage4_col7[1] <= stage3_col7[1];
                    stage4_col8[0] <= stage3_col8[0];
                    stage4_col8[1] <= stage3_col8[1];
                    stage4_col9[0] <= stage3_col9[0];
                    stage4_col9[1] <= stage3_col9[1];
                    stage4_col10[0] <= stage3_col10[0];
                    stage4_col10[1] <= stage3_col10[1];
                    stage4_col11[0] <= stage3_col11[0];
                    stage4_col11[1] <= stage3_col11[1];
                    stage4_col12[0] <= stage3_col12[0];
                    stage4_col12[1] <= stage3_col12[1];
                    stage4_col13[0] <= fa_s3_c13_n1_s;
                    stage4_col13[1] <= stage3_col13[3];
                    stage4_col14[0] <= fa_s3_c13_n1_c;
                    stage4_col14[1] <= fa_s3_c14_n2_s;
                    stage4_col15[0] <= fa_s3_c14_n2_c;
                    stage4_col15[1] <= fa_s3_c15_n3_s;
                    stage4_col16[0] <= fa_s3_c15_n3_c;
                    stage4_col16[1] <= fa_s3_c16_n4_s;
                    stage4_col17[0] <= fa_s3_c16_n4_c;
                    stage4_col17[1] <= fa_s3_c17_n5_s;
                    stage4_col18[0] <= fa_s3_c17_n5_c;
                    stage4_col18[1] <= fa_s3_c18_n6_s;
                    stage4_col19[0] <= fa_s3_c18_n6_c;
                    stage4_col19[1] <= fa_s3_c19_n7_s;
                    stage4_col19[2] <= stage3_col19[3];
                    stage4_col19[3] <= stage3_col19[4];
                    stage4_col20[0] <= fa_s3_c19_n7_c;
                    stage4_col20[1] <= fa_s3_c20_n8_s;
                    stage4_col20[2] <= stage3_col20[3];
                    stage4_col21[0] <= fa_s3_c20_n8_c;
                    stage4_col21[1] <= fa_s3_c21_n9_s;
                    stage4_col21[2] <= stage3_col21[3];
                    stage4_col22[0] <= fa_s3_c21_n9_c;
                    stage4_col22[1] <= fa_s3_c22_n10_s;
                    stage4_col22[2] <= stage3_col22[3];
                    stage4_col23[0] <= fa_s3_c22_n10_c;
                    stage4_col23[1] <= fa_s3_c23_n11_s;
                    stage4_col23[2] <= stage3_col23[3];
                    stage4_col24[0] <= fa_s3_c23_n11_c;
                    stage4_col24[1] <= fa_s3_c24_n12_s;
                    stage4_col24[2] <= stage3_col24[3];
                    stage4_col25[0] <= fa_s3_c24_n12_c;
                    stage4_col25[1] <= fa_s3_c25_n13_s;
                    stage4_col25[2] <= stage3_col25[3];
                    stage4_col26[0] <= fa_s3_c25_n13_c;
                    stage4_col26[1] <= fa_s3_c26_n14_s;
                    stage4_col26[2] <= stage3_col26[3];
                    stage4_col27[0] <= fa_s3_c26_n14_c;
                    stage4_col27[1] <= fa_s3_c27_n15_s;
                    stage4_col27[2] <= fa_s3_c27_n16_s;
                    stage4_col28[0] <= fa_s3_c27_n15_c;
                    stage4_col28[1] <= fa_s3_c27_n16_c;
                    stage4_col28[2] <= fa_s3_c28_n17_s;
                    stage4_col28[3] <= stage3_col28[3];
                    stage4_col28[4] <= stage3_col28[4];
                    stage4_col29[0] <= fa_s3_c28_n17_c;
                    stage4_col29[1] <= fa_s3_c29_n18_s;
                    stage4_col29[2] <= stage3_col29[3];
                    stage4_col29[3] <= stage3_col29[4];
                    stage4_col30[0] <= fa_s3_c29_n18_c;
                    stage4_col30[1] <= fa_s3_c30_n19_s;
                    stage4_col30[2] <= stage3_col30[3];
                    stage4_col30[3] <= stage3_col30[4];
                    stage4_col31[0] <= fa_s3_c30_n19_c;
                    stage4_col31[1] <= fa_s3_c31_n20_s;
                    stage4_col31[2] <= stage3_col31[3];
                    stage4_col31[3] <= stage3_col31[4];
                    stage4_col32[0] <= fa_s3_c31_n20_c;
                    stage4_col32[1] <= fa_s3_c32_n21_s;
                    stage4_col32[2] <= fa_s3_c32_n22_s;
                    stage4_col32[3] <= stage3_col32[6];
                    stage4_col33[0] <= fa_s3_c32_n21_c;
                    stage4_col33[1] <= fa_s3_c32_n22_c;
                    stage4_col33[2] <= fa_s3_c33_n23_s;
                    stage4_col33[3] <= fa_s3_c33_n24_s;
                    stage4_col34[0] <= fa_s3_c33_n23_c;
                    stage4_col34[1] <= fa_s3_c33_n24_c;
                    stage4_col34[2] <= fa_s3_c34_n25_s;
                    stage4_col34[3] <= fa_s3_c34_n26_s;
                    stage4_col35[0] <= fa_s3_c34_n25_c;
                    stage4_col35[1] <= fa_s3_c34_n26_c;
                    stage4_col35[2] <= fa_s3_c35_n27_s;
                    stage4_col35[3] <= fa_s3_c35_n28_s;
                    stage4_col36[0] <= fa_s3_c35_n27_c;
                    stage4_col36[1] <= fa_s3_c35_n28_c;
                    stage4_col36[2] <= fa_s3_c36_n29_s;
                    stage4_col36[3] <= fa_s3_c36_n30_s;
                    stage4_col37[0] <= fa_s3_c36_n29_c;
                    stage4_col37[1] <= fa_s3_c36_n30_c;
                    stage4_col37[2] <= fa_s3_c37_n31_s;
                    stage4_col37[3] <= fa_s3_c37_n32_s;
                    stage4_col38[0] <= fa_s3_c37_n31_c;
                    stage4_col38[1] <= fa_s3_c37_n32_c;
                    stage4_col38[2] <= fa_s3_c38_n33_s;
                    stage4_col38[3] <= fa_s3_c38_n34_s;
                    stage4_col39[0] <= fa_s3_c38_n33_c;
                    stage4_col39[1] <= fa_s3_c38_n34_c;
                    stage4_col39[2] <= fa_s3_c39_n35_s;
                    stage4_col39[3] <= fa_s3_c39_n36_s;
                    stage4_col40[0] <= fa_s3_c39_n35_c;
                    stage4_col40[1] <= fa_s3_c39_n36_c;
                    stage4_col40[2] <= fa_s3_c40_n37_s;
                    stage4_col40[3] <= fa_s3_c40_n38_s;
                    stage4_col40[4] <= stage3_col40[6];
                    stage4_col40[5] <= stage3_col40[7];
                    stage4_col41[0] <= fa_s3_c40_n37_c;
                    stage4_col41[1] <= fa_s3_c40_n38_c;
                    stage4_col41[2] <= fa_s3_c41_n39_s;
                    stage4_col41[3] <= fa_s3_c41_n40_s;
                    stage4_col41[4] <= stage3_col41[6];
                    stage4_col42[0] <= fa_s3_c41_n39_c;
                    stage4_col42[1] <= fa_s3_c41_n40_c;
                    stage4_col42[2] <= fa_s3_c42_n41_s;
                    stage4_col42[3] <= fa_s3_c42_n42_s;
                    stage4_col42[4] <= stage3_col42[6];
                    stage4_col43[0] <= fa_s3_c42_n41_c;
                    stage4_col43[1] <= fa_s3_c42_n42_c;
                    stage4_col43[2] <= fa_s3_c43_n43_s;
                    stage4_col43[3] <= fa_s3_c43_n44_s;
                    stage4_col43[4] <= stage3_col43[6];
                    stage4_col44[0] <= fa_s3_c43_n43_c;
                    stage4_col44[1] <= fa_s3_c43_n44_c;
                    stage4_col44[2] <= fa_s3_c44_n45_s;
                    stage4_col44[3] <= fa_s3_c44_n46_s;
                    stage4_col44[4] <= stage3_col44[6];
                    stage4_col45[0] <= fa_s3_c44_n45_c;
                    stage4_col45[1] <= fa_s3_c44_n46_c;
                    stage4_col45[2] <= fa_s3_c45_n47_s;
                    stage4_col45[3] <= fa_s3_c45_n48_s;
                    stage4_col45[4] <= stage3_col45[6];
                    stage4_col46[0] <= fa_s3_c45_n47_c;
                    stage4_col46[1] <= fa_s3_c45_n48_c;
                    stage4_col46[2] <= fa_s3_c46_n49_s;
                    stage4_col46[3] <= fa_s3_c46_n50_s;
                    stage4_col46[4] <= fa_s3_c46_n51_s;
                    stage4_col47[0] <= fa_s3_c46_n49_c;
                    stage4_col47[1] <= fa_s3_c46_n50_c;
                    stage4_col47[2] <= fa_s3_c46_n51_c;
                    stage4_col47[3] <= fa_s3_c47_n52_s;
                    stage4_col47[4] <= fa_s3_c47_n53_s;
                    stage4_col47[5] <= stage3_col47[6];
                    stage4_col47[6] <= stage3_col47[7];
                    stage4_col48[0] <= fa_s3_c47_n52_c;
                    stage4_col48[1] <= fa_s3_c47_n53_c;
                    stage4_col48[2] <= fa_s3_c48_n54_s;
                    stage4_col48[3] <= fa_s3_c48_n55_s;
                    stage4_col48[4] <= stage3_col48[6];
                    stage4_col48[5] <= stage3_col48[7];
                    stage4_col49[0] <= fa_s3_c48_n54_c;
                    stage4_col49[1] <= fa_s3_c48_n55_c;
                    stage4_col49[2] <= fa_s3_c49_n56_s;
                    stage4_col49[3] <= fa_s3_c49_n57_s;
                    stage4_col49[4] <= stage3_col49[6];
                    stage4_col49[5] <= stage3_col49[7];
                    stage4_col50[0] <= fa_s3_c49_n56_c;
                    stage4_col50[1] <= fa_s3_c49_n57_c;
                    stage4_col50[2] <= fa_s3_c50_n58_s;
                    stage4_col50[3] <= fa_s3_c50_n59_s;
                    stage4_col50[4] <= stage3_col50[6];
                    stage4_col50[5] <= stage3_col50[7];
                    stage4_col51[0] <= fa_s3_c50_n58_c;
                    stage4_col51[1] <= fa_s3_c50_n59_c;
                    stage4_col51[2] <= fa_s3_c51_n60_s;
                    stage4_col51[3] <= fa_s3_c51_n61_s;
                    stage4_col51[4] <= stage3_col51[6];
                    stage4_col51[5] <= stage3_col51[7];
                    stage4_col52[0] <= fa_s3_c51_n60_c;
                    stage4_col52[1] <= fa_s3_c51_n61_c;
                    stage4_col52[2] <= fa_s3_c52_n62_s;
                    stage4_col52[3] <= fa_s3_c52_n63_s;
                    stage4_col52[4] <= stage3_col52[6];
                    stage4_col52[5] <= stage3_col52[7];
                    stage4_col53[0] <= fa_s3_c52_n62_c;
                    stage4_col53[1] <= fa_s3_c52_n63_c;
                    stage4_col53[2] <= fa_s3_c53_n64_s;
                    stage4_col53[3] <= fa_s3_c53_n65_s;
                    stage4_col53[4] <= stage3_col53[6];
                    stage4_col53[5] <= stage3_col53[7];
                    stage4_col54[0] <= fa_s3_c53_n64_c;
                    stage4_col54[1] <= fa_s3_c53_n65_c;
                    stage4_col54[2] <= fa_s3_c54_n66_s;
                    stage4_col54[3] <= fa_s3_c54_n67_s;
                    stage4_col54[4] <= fa_s3_c54_n68_s;
                    stage4_col54[5] <= stage3_col54[9];
                    stage4_col55[0] <= fa_s3_c54_n66_c;
                    stage4_col55[1] <= fa_s3_c54_n67_c;
                    stage4_col55[2] <= fa_s3_c54_n68_c;
                    stage4_col55[3] <= fa_s3_c55_n69_s;
                    stage4_col55[4] <= fa_s3_c55_n70_s;
                    stage4_col55[5] <= fa_s3_c55_n71_s;
                    stage4_col56[0] <= fa_s3_c55_n69_c;
                    stage4_col56[1] <= fa_s3_c55_n70_c;
                    stage4_col56[2] <= fa_s3_c55_n71_c;
                    stage4_col56[3] <= fa_s3_c56_n72_s;
                    stage4_col56[4] <= fa_s3_c56_n73_s;
                    stage4_col56[5] <= fa_s3_c56_n74_s;
                    stage4_col57[0] <= fa_s3_c56_n72_c;
                    stage4_col57[1] <= fa_s3_c56_n73_c;
                    stage4_col57[2] <= fa_s3_c56_n74_c;
                    stage4_col57[3] <= fa_s3_c57_n75_s;
                    stage4_col57[4] <= fa_s3_c57_n76_s;
                    stage4_col57[5] <= fa_s3_c57_n77_s;
                    stage4_col58[0] <= fa_s3_c57_n75_c;
                    stage4_col58[1] <= fa_s3_c57_n76_c;
                    stage4_col58[2] <= fa_s3_c57_n77_c;
                    stage4_col58[3] <= fa_s3_c58_n78_s;
                    stage4_col58[4] <= fa_s3_c58_n79_s;
                    stage4_col58[5] <= fa_s3_c58_n80_s;
                    stage4_col59[0] <= fa_s3_c58_n78_c;
                    stage4_col59[1] <= fa_s3_c58_n79_c;
                    stage4_col59[2] <= fa_s3_c58_n80_c;
                    stage4_col59[3] <= fa_s3_c59_n81_s;
                    stage4_col59[4] <= fa_s3_c59_n82_s;
                    stage4_col59[5] <= fa_s3_c59_n83_s;
                    stage4_col59[6] <= stage3_col59[9];
                    stage4_col59[7] <= stage3_col59[10];
                    stage4_col60[0] <= fa_s3_c59_n81_c;
                    stage4_col60[1] <= fa_s3_c59_n82_c;
                    stage4_col60[2] <= fa_s3_c59_n83_c;
                    stage4_col60[3] <= fa_s3_c60_n84_s;
                    stage4_col60[4] <= fa_s3_c60_n85_s;
                    stage4_col60[5] <= fa_s3_c60_n86_s;
                    stage4_col60[6] <= stage3_col60[9];
                    stage4_col61[0] <= fa_s3_c60_n84_c;
                    stage4_col61[1] <= fa_s3_c60_n85_c;
                    stage4_col61[2] <= fa_s3_c60_n86_c;
                    stage4_col61[3] <= fa_s3_c61_n87_s;
                    stage4_col61[4] <= fa_s3_c61_n88_s;
                    stage4_col61[5] <= fa_s3_c61_n89_s;
                    stage4_col61[6] <= stage3_col61[9];
                    stage4_col62[0] <= fa_s3_c61_n87_c;
                    stage4_col62[1] <= fa_s3_c61_n88_c;
                    stage4_col62[2] <= fa_s3_c61_n89_c;
                    stage4_col62[3] <= fa_s3_c62_n90_s;
                    stage4_col62[4] <= fa_s3_c62_n91_s;
                    stage4_col62[5] <= fa_s3_c62_n92_s;
                    stage4_col62[6] <= stage3_col62[9];
                    stage4_col63[0] <= fa_s3_c62_n90_c;
                    stage4_col63[1] <= fa_s3_c62_n91_c;
                    stage4_col63[2] <= fa_s3_c62_n92_c;
                    stage4_col63[3] <= fa_s3_c63_n93_s;
                    stage4_col63[4] <= fa_s3_c63_n94_s;
                    stage4_col63[5] <= fa_s3_c63_n95_s;
                    stage4_col63[6] <= stage3_col63[9];
                    stage4_col64[0] <= fa_s3_c63_n93_c;
                    stage4_col64[1] <= fa_s3_c63_n94_c;
                    stage4_col64[2] <= fa_s3_c63_n95_c;
                    stage4_col64[3] <= fa_s3_c64_n96_s;
                    stage4_col64[4] <= fa_s3_c64_n97_s;
                    stage4_col64[5] <= fa_s3_c64_n98_s;
                    stage4_col64[6] <= stage3_col64[9];
                    stage4_col64[7] <= stage3_col64[10];
                    stage4_col65[0] <= fa_s3_c64_n96_c;
                    stage4_col65[1] <= fa_s3_c64_n97_c;
                    stage4_col65[2] <= fa_s3_c64_n98_c;
                    stage4_col65[3] <= fa_s3_c65_n99_s;
                    stage4_col65[4] <= fa_s3_c65_n100_s;
                    stage4_col65[5] <= fa_s3_c65_n101_s;
                    stage4_col65[6] <= stage3_col65[9];
                    stage4_col66[0] <= fa_s3_c65_n99_c;
                    stage4_col66[1] <= fa_s3_c65_n100_c;
                    stage4_col66[2] <= fa_s3_c65_n101_c;
                    stage4_col66[3] <= fa_s3_c66_n102_s;
                    stage4_col66[4] <= fa_s3_c66_n103_s;
                    stage4_col66[5] <= fa_s3_c66_n104_s;
                    stage4_col66[6] <= stage3_col66[9];
                    stage4_col66[7] <= stage3_col66[10];
                    stage4_col67[0] <= fa_s3_c66_n102_c;
                    stage4_col67[1] <= fa_s3_c66_n103_c;
                    stage4_col67[2] <= fa_s3_c66_n104_c;
                    stage4_col67[3] <= fa_s3_c67_n105_s;
                    stage4_col67[4] <= fa_s3_c67_n106_s;
                    stage4_col67[5] <= fa_s3_c67_n107_s;
                    stage4_col67[6] <= stage3_col67[9];
                    stage4_col68[0] <= fa_s3_c67_n105_c;
                    stage4_col68[1] <= fa_s3_c67_n106_c;
                    stage4_col68[2] <= fa_s3_c67_n107_c;
                    stage4_col68[3] <= fa_s3_c68_n108_s;
                    stage4_col68[4] <= fa_s3_c68_n109_s;
                    stage4_col68[5] <= fa_s3_c68_n110_s;
                    stage4_col68[6] <= stage3_col68[9];
                    stage4_col68[7] <= stage3_col68[10];
                    stage4_col69[0] <= fa_s3_c68_n108_c;
                    stage4_col69[1] <= fa_s3_c68_n109_c;
                    stage4_col69[2] <= fa_s3_c68_n110_c;
                    stage4_col69[3] <= fa_s3_c69_n111_s;
                    stage4_col69[4] <= fa_s3_c69_n112_s;
                    stage4_col69[5] <= fa_s3_c69_n113_s;
                    stage4_col69[6] <= stage3_col69[9];
                    stage4_col70[0] <= fa_s3_c69_n111_c;
                    stage4_col70[1] <= fa_s3_c69_n112_c;
                    stage4_col70[2] <= fa_s3_c69_n113_c;
                    stage4_col70[3] <= fa_s3_c70_n114_s;
                    stage4_col70[4] <= fa_s3_c70_n115_s;
                    stage4_col70[5] <= fa_s3_c70_n116_s;
                    stage4_col70[6] <= stage3_col70[9];
                    stage4_col70[7] <= stage3_col70[10];
                    stage4_col71[0] <= fa_s3_c70_n114_c;
                    stage4_col71[1] <= fa_s3_c70_n115_c;
                    stage4_col71[2] <= fa_s3_c70_n116_c;
                    stage4_col71[3] <= fa_s3_c71_n117_s;
                    stage4_col71[4] <= fa_s3_c71_n118_s;
                    stage4_col71[5] <= fa_s3_c71_n119_s;
                    stage4_col71[6] <= stage3_col71[9];
                    stage4_col72[0] <= fa_s3_c71_n117_c;
                    stage4_col72[1] <= fa_s3_c71_n118_c;
                    stage4_col72[2] <= fa_s3_c71_n119_c;
                    stage4_col72[3] <= fa_s3_c72_n120_s;
                    stage4_col72[4] <= fa_s3_c72_n121_s;
                    stage4_col72[5] <= fa_s3_c72_n122_s;
                    stage4_col72[6] <= stage3_col72[9];
                    stage4_col72[7] <= stage3_col72[10];
                    stage4_col73[0] <= fa_s3_c72_n120_c;
                    stage4_col73[1] <= fa_s3_c72_n121_c;
                    stage4_col73[2] <= fa_s3_c72_n122_c;
                    stage4_col73[3] <= fa_s3_c73_n123_s;
                    stage4_col73[4] <= fa_s3_c73_n124_s;
                    stage4_col73[5] <= fa_s3_c73_n125_s;
                    stage4_col73[6] <= stage3_col73[9];
                    stage4_col74[0] <= fa_s3_c73_n123_c;
                    stage4_col74[1] <= fa_s3_c73_n124_c;
                    stage4_col74[2] <= fa_s3_c73_n125_c;
                    stage4_col74[3] <= fa_s3_c74_n126_s;
                    stage4_col74[4] <= fa_s3_c74_n127_s;
                    stage4_col74[5] <= fa_s3_c74_n128_s;
                    stage4_col74[6] <= stage3_col74[9];
                    stage4_col74[7] <= stage3_col74[10];
                    stage4_col75[0] <= fa_s3_c74_n126_c;
                    stage4_col75[1] <= fa_s3_c74_n127_c;
                    stage4_col75[2] <= fa_s3_c74_n128_c;
                    stage4_col75[3] <= fa_s3_c75_n129_s;
                    stage4_col75[4] <= fa_s3_c75_n130_s;
                    stage4_col75[5] <= fa_s3_c75_n131_s;
                    stage4_col75[6] <= stage3_col75[9];
                    stage4_col76[0] <= fa_s3_c75_n129_c;
                    stage4_col76[1] <= fa_s3_c75_n130_c;
                    stage4_col76[2] <= fa_s3_c75_n131_c;
                    stage4_col76[3] <= fa_s3_c76_n132_s;
                    stage4_col76[4] <= fa_s3_c76_n133_s;
                    stage4_col76[5] <= fa_s3_c76_n134_s;
                    stage4_col76[6] <= stage3_col76[9];
                    stage4_col76[7] <= stage3_col76[10];
                    stage4_col77[0] <= fa_s3_c76_n132_c;
                    stage4_col77[1] <= fa_s3_c76_n133_c;
                    stage4_col77[2] <= fa_s3_c76_n134_c;
                    stage4_col77[3] <= fa_s3_c77_n135_s;
                    stage4_col77[4] <= fa_s3_c77_n136_s;
                    stage4_col77[5] <= fa_s3_c77_n137_s;
                    stage4_col77[6] <= stage3_col77[9];
                    stage4_col78[0] <= fa_s3_c77_n135_c;
                    stage4_col78[1] <= fa_s3_c77_n136_c;
                    stage4_col78[2] <= fa_s3_c77_n137_c;
                    stage4_col78[3] <= fa_s3_c78_n138_s;
                    stage4_col78[4] <= fa_s3_c78_n139_s;
                    stage4_col78[5] <= fa_s3_c78_n140_s;
                    stage4_col78[6] <= stage3_col78[9];
                    stage4_col78[7] <= stage3_col78[10];
                    stage4_col79[0] <= fa_s3_c78_n138_c;
                    stage4_col79[1] <= fa_s3_c78_n139_c;
                    stage4_col79[2] <= fa_s3_c78_n140_c;
                    stage4_col79[3] <= fa_s3_c79_n141_s;
                    stage4_col79[4] <= fa_s3_c79_n142_s;
                    stage4_col79[5] <= fa_s3_c79_n143_s;
                    stage4_col79[6] <= stage3_col79[9];
                    stage4_col80[0] <= fa_s3_c79_n141_c;
                    stage4_col80[1] <= fa_s3_c79_n142_c;
                    stage4_col80[2] <= fa_s3_c79_n143_c;
                    stage4_col80[3] <= fa_s3_c80_n144_s;
                    stage4_col80[4] <= fa_s3_c80_n145_s;
                    stage4_col80[5] <= fa_s3_c80_n146_s;
                    stage4_col80[6] <= stage3_col80[9];
                    stage4_col80[7] <= stage3_col80[10];
                    stage4_col81[0] <= fa_s3_c80_n144_c;
                    stage4_col81[1] <= fa_s3_c80_n145_c;
                    stage4_col81[2] <= fa_s3_c80_n146_c;
                    stage4_col81[3] <= fa_s3_c81_n147_s;
                    stage4_col81[4] <= fa_s3_c81_n148_s;
                    stage4_col81[5] <= fa_s3_c81_n149_s;
                    stage4_col81[6] <= stage3_col81[9];
                    stage4_col82[0] <= fa_s3_c81_n147_c;
                    stage4_col82[1] <= fa_s3_c81_n148_c;
                    stage4_col82[2] <= fa_s3_c81_n149_c;
                    stage4_col82[3] <= fa_s3_c82_n150_s;
                    stage4_col82[4] <= fa_s3_c82_n151_s;
                    stage4_col82[5] <= fa_s3_c82_n152_s;
                    stage4_col82[6] <= stage3_col82[9];
                    stage4_col82[7] <= stage3_col82[10];
                    stage4_col83[0] <= fa_s3_c82_n150_c;
                    stage4_col83[1] <= fa_s3_c82_n151_c;
                    stage4_col83[2] <= fa_s3_c82_n152_c;
                    stage4_col83[3] <= fa_s3_c83_n153_s;
                    stage4_col83[4] <= fa_s3_c83_n154_s;
                    stage4_col83[5] <= fa_s3_c83_n155_s;
                    stage4_col83[6] <= stage3_col83[9];
                    stage4_col84[0] <= fa_s3_c83_n153_c;
                    stage4_col84[1] <= fa_s3_c83_n154_c;
                    stage4_col84[2] <= fa_s3_c83_n155_c;
                    stage4_col84[3] <= fa_s3_c84_n156_s;
                    stage4_col84[4] <= fa_s3_c84_n157_s;
                    stage4_col84[5] <= fa_s3_c84_n158_s;
                    stage4_col84[6] <= stage3_col84[9];
                    stage4_col84[7] <= stage3_col84[10];
                    stage4_col85[0] <= fa_s3_c84_n156_c;
                    stage4_col85[1] <= fa_s3_c84_n157_c;
                    stage4_col85[2] <= fa_s3_c84_n158_c;
                    stage4_col85[3] <= fa_s3_c85_n159_s;
                    stage4_col85[4] <= fa_s3_c85_n160_s;
                    stage4_col85[5] <= fa_s3_c85_n161_s;
                    stage4_col85[6] <= stage3_col85[9];
                    stage4_col86[0] <= fa_s3_c85_n159_c;
                    stage4_col86[1] <= fa_s3_c85_n160_c;
                    stage4_col86[2] <= fa_s3_c85_n161_c;
                    stage4_col86[3] <= fa_s3_c86_n162_s;
                    stage4_col86[4] <= fa_s3_c86_n163_s;
                    stage4_col86[5] <= fa_s3_c86_n164_s;
                    stage4_col86[6] <= stage3_col86[9];
                    stage4_col86[7] <= stage3_col86[10];
                    stage4_col87[0] <= fa_s3_c86_n162_c;
                    stage4_col87[1] <= fa_s3_c86_n163_c;
                    stage4_col87[2] <= fa_s3_c86_n164_c;
                    stage4_col87[3] <= fa_s3_c87_n165_s;
                    stage4_col87[4] <= fa_s3_c87_n166_s;
                    stage4_col87[5] <= fa_s3_c87_n167_s;
                    stage4_col87[6] <= stage3_col87[9];
                    stage4_col88[0] <= fa_s3_c87_n165_c;
                    stage4_col88[1] <= fa_s3_c87_n166_c;
                    stage4_col88[2] <= fa_s3_c87_n167_c;
                    stage4_col88[3] <= fa_s3_c88_n168_s;
                    stage4_col88[4] <= fa_s3_c88_n169_s;
                    stage4_col88[5] <= fa_s3_c88_n170_s;
                    stage4_col88[6] <= stage3_col88[9];
                    stage4_col88[7] <= stage3_col88[10];
                    stage4_col89[0] <= fa_s3_c88_n168_c;
                    stage4_col89[1] <= fa_s3_c88_n169_c;
                    stage4_col89[2] <= fa_s3_c88_n170_c;
                    stage4_col89[3] <= fa_s3_c89_n171_s;
                    stage4_col89[4] <= fa_s3_c89_n172_s;
                    stage4_col89[5] <= fa_s3_c89_n173_s;
                    stage4_col89[6] <= stage3_col89[9];
                    stage4_col90[0] <= fa_s3_c89_n171_c;
                    stage4_col90[1] <= fa_s3_c89_n172_c;
                    stage4_col90[2] <= fa_s3_c89_n173_c;
                    stage4_col90[3] <= fa_s3_c90_n174_s;
                    stage4_col90[4] <= fa_s3_c90_n175_s;
                    stage4_col90[5] <= fa_s3_c90_n176_s;
                    stage4_col90[6] <= stage3_col90[9];
                    stage4_col90[7] <= stage3_col90[10];
                    stage4_col91[0] <= fa_s3_c90_n174_c;
                    stage4_col91[1] <= fa_s3_c90_n175_c;
                    stage4_col91[2] <= fa_s3_c90_n176_c;
                    stage4_col91[3] <= fa_s3_c91_n177_s;
                    stage4_col91[4] <= fa_s3_c91_n178_s;
                    stage4_col91[5] <= fa_s3_c91_n179_s;
                    stage4_col91[6] <= stage3_col91[9];
                    stage4_col92[0] <= fa_s3_c91_n177_c;
                    stage4_col92[1] <= fa_s3_c91_n178_c;
                    stage4_col92[2] <= fa_s3_c91_n179_c;
                    stage4_col92[3] <= fa_s3_c92_n180_s;
                    stage4_col92[4] <= fa_s3_c92_n181_s;
                    stage4_col92[5] <= fa_s3_c92_n182_s;
                    stage4_col92[6] <= stage3_col92[9];
                    stage4_col92[7] <= stage3_col92[10];
                    stage4_col93[0] <= fa_s3_c92_n180_c;
                    stage4_col93[1] <= fa_s3_c92_n181_c;
                    stage4_col93[2] <= fa_s3_c92_n182_c;
                    stage4_col93[3] <= fa_s3_c93_n183_s;
                    stage4_col93[4] <= fa_s3_c93_n184_s;
                    stage4_col93[5] <= fa_s3_c93_n185_s;
                    stage4_col93[6] <= stage3_col93[9];
                    stage4_col94[0] <= fa_s3_c93_n183_c;
                    stage4_col94[1] <= fa_s3_c93_n184_c;
                    stage4_col94[2] <= fa_s3_c93_n185_c;
                    stage4_col94[3] <= fa_s3_c94_n186_s;
                    stage4_col94[4] <= fa_s3_c94_n187_s;
                    stage4_col94[5] <= fa_s3_c94_n188_s;
                    stage4_col94[6] <= stage3_col94[9];
                    stage4_col94[7] <= stage3_col94[10];
                    stage4_col95[0] <= fa_s3_c94_n186_c;
                    stage4_col95[1] <= fa_s3_c94_n187_c;
                    stage4_col95[2] <= fa_s3_c94_n188_c;
                    stage4_col95[3] <= fa_s3_c95_n189_s;
                    stage4_col95[4] <= fa_s3_c95_n190_s;
                    stage4_col95[5] <= fa_s3_c95_n191_s;
                    stage4_col95[6] <= stage3_col95[9];
                    stage4_col96[0] <= fa_s3_c95_n189_c;
                    stage4_col96[1] <= fa_s3_c95_n190_c;
                    stage4_col96[2] <= fa_s3_c95_n191_c;
                    stage4_col96[3] <= fa_s3_c96_n192_s;
                    stage4_col96[4] <= fa_s3_c96_n193_s;
                    stage4_col96[5] <= fa_s3_c96_n194_s;
                    stage4_col96[6] <= stage3_col96[9];
                    stage4_col96[7] <= stage3_col96[10];
                    stage4_col97[0] <= fa_s3_c96_n192_c;
                    stage4_col97[1] <= fa_s3_c96_n193_c;
                    stage4_col97[2] <= fa_s3_c96_n194_c;
                    stage4_col97[3] <= fa_s3_c97_n195_s;
                    stage4_col97[4] <= fa_s3_c97_n196_s;
                    stage4_col97[5] <= fa_s3_c97_n197_s;
                    stage4_col97[6] <= stage3_col97[9];
                    stage4_col98[0] <= fa_s3_c97_n195_c;
                    stage4_col98[1] <= fa_s3_c97_n196_c;
                    stage4_col98[2] <= fa_s3_c97_n197_c;
                    stage4_col98[3] <= fa_s3_c98_n198_s;
                    stage4_col98[4] <= fa_s3_c98_n199_s;
                    stage4_col98[5] <= fa_s3_c98_n200_s;
                    stage4_col98[6] <= stage3_col98[9];
                    stage4_col98[7] <= stage3_col98[10];
                    stage4_col99[0] <= fa_s3_c98_n198_c;
                    stage4_col99[1] <= fa_s3_c98_n199_c;
                    stage4_col99[2] <= fa_s3_c98_n200_c;
                    stage4_col99[3] <= fa_s3_c99_n201_s;
                    stage4_col99[4] <= fa_s3_c99_n202_s;
                    stage4_col99[5] <= fa_s3_c99_n203_s;
                    stage4_col99[6] <= stage3_col99[9];
                    stage4_col100[0] <= fa_s3_c99_n201_c;
                    stage4_col100[1] <= fa_s3_c99_n202_c;
                    stage4_col100[2] <= fa_s3_c99_n203_c;
                    stage4_col100[3] <= fa_s3_c100_n204_s;
                    stage4_col100[4] <= fa_s3_c100_n205_s;
                    stage4_col100[5] <= fa_s3_c100_n206_s;
                    stage4_col100[6] <= stage3_col100[9];
                    stage4_col100[7] <= stage3_col100[10];
                    stage4_col101[0] <= fa_s3_c100_n204_c;
                    stage4_col101[1] <= fa_s3_c100_n205_c;
                    stage4_col101[2] <= fa_s3_c100_n206_c;
                    stage4_col101[3] <= fa_s3_c101_n207_s;
                    stage4_col101[4] <= fa_s3_c101_n208_s;
                    stage4_col101[5] <= fa_s3_c101_n209_s;
                    stage4_col101[6] <= stage3_col101[9];
                    stage4_col102[0] <= fa_s3_c101_n207_c;
                    stage4_col102[1] <= fa_s3_c101_n208_c;
                    stage4_col102[2] <= fa_s3_c101_n209_c;
                    stage4_col102[3] <= fa_s3_c102_n210_s;
                    stage4_col102[4] <= fa_s3_c102_n211_s;
                    stage4_col102[5] <= fa_s3_c102_n212_s;
                    stage4_col102[6] <= stage3_col102[9];
                    stage4_col102[7] <= stage3_col102[10];
                    stage4_col103[0] <= fa_s3_c102_n210_c;
                    stage4_col103[1] <= fa_s3_c102_n211_c;
                    stage4_col103[2] <= fa_s3_c102_n212_c;
                    stage4_col103[3] <= fa_s3_c103_n213_s;
                    stage4_col103[4] <= fa_s3_c103_n214_s;
                    stage4_col103[5] <= fa_s3_c103_n215_s;
                    stage4_col103[6] <= stage3_col103[9];
                    stage4_col104[0] <= fa_s3_c103_n213_c;
                    stage4_col104[1] <= fa_s3_c103_n214_c;
                    stage4_col104[2] <= fa_s3_c103_n215_c;
                    stage4_col104[3] <= fa_s3_c104_n216_s;
                    stage4_col104[4] <= fa_s3_c104_n217_s;
                    stage4_col104[5] <= fa_s3_c104_n218_s;
                    stage4_col104[6] <= stage3_col104[9];
                    stage4_col104[7] <= stage3_col104[10];
                    stage4_col105[0] <= fa_s3_c104_n216_c;
                    stage4_col105[1] <= fa_s3_c104_n217_c;
                    stage4_col105[2] <= fa_s3_c104_n218_c;
                    stage4_col105[3] <= fa_s3_c105_n219_s;
                    stage4_col105[4] <= fa_s3_c105_n220_s;
                    stage4_col105[5] <= fa_s3_c105_n221_s;
                    stage4_col105[6] <= stage3_col105[9];
                    stage4_col106[0] <= fa_s3_c105_n219_c;
                    stage4_col106[1] <= fa_s3_c105_n220_c;
                    stage4_col106[2] <= fa_s3_c105_n221_c;
                    stage4_col106[3] <= fa_s3_c106_n222_s;
                    stage4_col106[4] <= fa_s3_c106_n223_s;
                    stage4_col106[5] <= fa_s3_c106_n224_s;
                    stage4_col106[6] <= stage3_col106[9];
                    stage4_col106[7] <= stage3_col106[10];
                    stage4_col107[0] <= fa_s3_c106_n222_c;
                    stage4_col107[1] <= fa_s3_c106_n223_c;
                    stage4_col107[2] <= fa_s3_c106_n224_c;
                    stage4_col107[3] <= fa_s3_c107_n225_s;
                    stage4_col107[4] <= fa_s3_c107_n226_s;
                    stage4_col107[5] <= fa_s3_c107_n227_s;
                    stage4_col107[6] <= stage3_col107[9];
                    stage4_col108[0] <= fa_s3_c107_n225_c;
                    stage4_col108[1] <= fa_s3_c107_n226_c;
                    stage4_col108[2] <= fa_s3_c107_n227_c;
                    stage4_col108[3] <= fa_s3_c108_n228_s;
                    stage4_col108[4] <= fa_s3_c108_n229_s;
                    stage4_col108[5] <= fa_s3_c108_n230_s;
                    stage4_col108[6] <= stage3_col108[9];
                    stage4_col108[7] <= stage3_col108[10];
                    stage4_col109[0] <= fa_s3_c108_n228_c;
                    stage4_col109[1] <= fa_s3_c108_n229_c;
                    stage4_col109[2] <= fa_s3_c108_n230_c;
                    stage4_col109[3] <= fa_s3_c109_n231_s;
                    stage4_col109[4] <= fa_s3_c109_n232_s;
                    stage4_col109[5] <= fa_s3_c109_n233_s;
                    stage4_col109[6] <= stage3_col109[9];
                    stage4_col110[0] <= fa_s3_c109_n231_c;
                    stage4_col110[1] <= fa_s3_c109_n232_c;
                    stage4_col110[2] <= fa_s3_c109_n233_c;
                    stage4_col110[3] <= fa_s3_c110_n234_s;
                    stage4_col110[4] <= fa_s3_c110_n235_s;
                    stage4_col110[5] <= fa_s3_c110_n236_s;
                    stage4_col110[6] <= stage3_col110[9];
                    stage4_col110[7] <= stage3_col110[10];
                    stage4_col111[0] <= fa_s3_c110_n234_c;
                    stage4_col111[1] <= fa_s3_c110_n235_c;
                    stage4_col111[2] <= fa_s3_c110_n236_c;
                    stage4_col111[3] <= fa_s3_c111_n237_s;
                    stage4_col111[4] <= fa_s3_c111_n238_s;
                    stage4_col111[5] <= fa_s3_c111_n239_s;
                    stage4_col111[6] <= stage3_col111[9];
                    stage4_col112[0] <= fa_s3_c111_n237_c;
                    stage4_col112[1] <= fa_s3_c111_n238_c;
                    stage4_col112[2] <= fa_s3_c111_n239_c;
                    stage4_col112[3] <= fa_s3_c112_n240_s;
                    stage4_col112[4] <= fa_s3_c112_n241_s;
                    stage4_col112[5] <= fa_s3_c112_n242_s;
                    stage4_col112[6] <= stage3_col112[9];
                    stage4_col112[7] <= stage3_col112[10];
                    stage4_col113[0] <= fa_s3_c112_n240_c;
                    stage4_col113[1] <= fa_s3_c112_n241_c;
                    stage4_col113[2] <= fa_s3_c112_n242_c;
                    stage4_col113[3] <= fa_s3_c113_n243_s;
                    stage4_col113[4] <= fa_s3_c113_n244_s;
                    stage4_col113[5] <= fa_s3_c113_n245_s;
                    stage4_col113[6] <= stage3_col113[9];
                    stage4_col114[0] <= fa_s3_c113_n243_c;
                    stage4_col114[1] <= fa_s3_c113_n244_c;
                    stage4_col114[2] <= fa_s3_c113_n245_c;
                    stage4_col114[3] <= fa_s3_c114_n246_s;
                    stage4_col114[4] <= fa_s3_c114_n247_s;
                    stage4_col114[5] <= fa_s3_c114_n248_s;
                    stage4_col114[6] <= stage3_col114[9];
                    stage4_col114[7] <= stage3_col114[10];
                    stage4_col115[0] <= fa_s3_c114_n246_c;
                    stage4_col115[1] <= fa_s3_c114_n247_c;
                    stage4_col115[2] <= fa_s3_c114_n248_c;
                    stage4_col115[3] <= fa_s3_c115_n249_s;
                    stage4_col115[4] <= fa_s3_c115_n250_s;
                    stage4_col115[5] <= fa_s3_c115_n251_s;
                    stage4_col115[6] <= stage3_col115[9];
                    stage4_col116[0] <= fa_s3_c115_n249_c;
                    stage4_col116[1] <= fa_s3_c115_n250_c;
                    stage4_col116[2] <= fa_s3_c115_n251_c;
                    stage4_col116[3] <= fa_s3_c116_n252_s;
                    stage4_col116[4] <= fa_s3_c116_n253_s;
                    stage4_col116[5] <= fa_s3_c116_n254_s;
                    stage4_col116[6] <= stage3_col116[9];
                    stage4_col116[7] <= stage3_col116[10];
                    stage4_col117[0] <= fa_s3_c116_n252_c;
                    stage4_col117[1] <= fa_s3_c116_n253_c;
                    stage4_col117[2] <= fa_s3_c116_n254_c;
                    stage4_col117[3] <= fa_s3_c117_n255_s;
                    stage4_col117[4] <= fa_s3_c117_n256_s;
                    stage4_col117[5] <= fa_s3_c117_n257_s;
                    stage4_col117[6] <= stage3_col117[9];
                    stage4_col118[0] <= fa_s3_c117_n255_c;
                    stage4_col118[1] <= fa_s3_c117_n256_c;
                    stage4_col118[2] <= fa_s3_c117_n257_c;
                    stage4_col118[3] <= fa_s3_c118_n258_s;
                    stage4_col118[4] <= fa_s3_c118_n259_s;
                    stage4_col118[5] <= fa_s3_c118_n260_s;
                    stage4_col118[6] <= stage3_col118[9];
                    stage4_col118[7] <= stage3_col118[10];
                    stage4_col119[0] <= fa_s3_c118_n258_c;
                    stage4_col119[1] <= fa_s3_c118_n259_c;
                    stage4_col119[2] <= fa_s3_c118_n260_c;
                    stage4_col119[3] <= fa_s3_c119_n261_s;
                    stage4_col119[4] <= fa_s3_c119_n262_s;
                    stage4_col119[5] <= fa_s3_c119_n263_s;
                    stage4_col119[6] <= stage3_col119[9];
                    stage4_col120[0] <= fa_s3_c119_n261_c;
                    stage4_col120[1] <= fa_s3_c119_n262_c;
                    stage4_col120[2] <= fa_s3_c119_n263_c;
                    stage4_col120[3] <= fa_s3_c120_n264_s;
                    stage4_col120[4] <= fa_s3_c120_n265_s;
                    stage4_col120[5] <= fa_s3_c120_n266_s;
                    stage4_col120[6] <= stage3_col120[9];
                    stage4_col120[7] <= stage3_col120[10];
                    stage4_col121[0] <= fa_s3_c120_n264_c;
                    stage4_col121[1] <= fa_s3_c120_n265_c;
                    stage4_col121[2] <= fa_s3_c120_n266_c;
                    stage4_col121[3] <= fa_s3_c121_n267_s;
                    stage4_col121[4] <= fa_s3_c121_n268_s;
                    stage4_col121[5] <= fa_s3_c121_n269_s;
                    stage4_col121[6] <= stage3_col121[9];
                    stage4_col122[0] <= fa_s3_c121_n267_c;
                    stage4_col122[1] <= fa_s3_c121_n268_c;
                    stage4_col122[2] <= fa_s3_c121_n269_c;
                    stage4_col122[3] <= fa_s3_c122_n270_s;
                    stage4_col122[4] <= fa_s3_c122_n271_s;
                    stage4_col122[5] <= fa_s3_c122_n272_s;
                    stage4_col122[6] <= stage3_col122[9];
                    stage4_col122[7] <= stage3_col122[10];
                    stage4_col123[0] <= fa_s3_c122_n270_c;
                    stage4_col123[1] <= fa_s3_c122_n271_c;
                    stage4_col123[2] <= fa_s3_c122_n272_c;
                    stage4_col123[3] <= fa_s3_c123_n273_s;
                    stage4_col123[4] <= fa_s3_c123_n274_s;
                    stage4_col123[5] <= fa_s3_c123_n275_s;
                    stage4_col123[6] <= stage3_col123[9];
                    stage4_col124[0] <= fa_s3_c123_n273_c;
                    stage4_col124[1] <= fa_s3_c123_n274_c;
                    stage4_col124[2] <= fa_s3_c123_n275_c;
                    stage4_col124[3] <= fa_s3_c124_n276_s;
                    stage4_col124[4] <= fa_s3_c124_n277_s;
                    stage4_col124[5] <= fa_s3_c124_n278_s;
                    stage4_col124[6] <= stage3_col124[9];
                    stage4_col124[7] <= stage3_col124[10];
                    stage4_col125[0] <= fa_s3_c124_n276_c;
                    stage4_col125[1] <= fa_s3_c124_n277_c;
                    stage4_col125[2] <= fa_s3_c124_n278_c;
                    stage4_col125[3] <= fa_s3_c125_n279_s;
                    stage4_col125[4] <= fa_s3_c125_n280_s;
                    stage4_col125[5] <= fa_s3_c125_n281_s;
                    stage4_col125[6] <= stage3_col125[9];
                    stage4_col126[0] <= fa_s3_c125_n279_c;
                    stage4_col126[1] <= fa_s3_c125_n280_c;
                    stage4_col126[2] <= fa_s3_c125_n281_c;
                    stage4_col126[3] <= fa_s3_c126_n282_s;
                    stage4_col126[4] <= fa_s3_c126_n283_s;
                    stage4_col126[5] <= fa_s3_c126_n284_s;
                    stage4_col126[6] <= stage3_col126[9];
                    stage4_col126[7] <= stage3_col126[10];
                    stage4_col127[0] <= fa_s3_c126_n282_c;
                    stage4_col127[1] <= fa_s3_c126_n283_c;
                    stage4_col127[2] <= fa_s3_c126_n284_c;
                    stage4_col127[3] <= stage3_col127[0];
                    stage4_col127[4] <= stage3_col127[1];
                    stage4_col127[5] <= stage3_col127[2];
                    stage4_col127[6] <= stage3_col127[3];
                    stage4_col127[7] <= stage3_col127[4];
                    stage4_col127[8] <= stage3_col127[5];
                    stage4_col127[9] <= stage3_col127[6];
                    stage4_col127[10] <= stage3_col127[7];
                    stage4_col127[11] <= stage3_col127[8];
                    stage4_col127[12] <= stage3_col127[9];
                    stage4_col127[13] <= stage3_col127[10];
                    stage4_col127[14] <= stage3_col127[11];
                    stage4_col127[15] <= stage3_col127[12];
                    stage4_col127[16] <= stage3_col127[13];
                    stage4_col127[17] <= stage3_col127[14];
                    stage4_col127[18] <= stage3_col127[15];
                    stage4_col127[19] <= stage3_col127[16];
                    stage4_col127[20] <= stage3_col127[17];
                    stage4_col127[21] <= stage3_col127[18];
                    stage4_col127[22] <= stage3_col127[19];
                    stage4_col127[23] <= stage3_col127[20];
                    stage4_col127[24] <= stage3_col127[21];
                    stage4_col127[25] <= stage3_col127[22];
                    stage4_col127[26] <= stage3_col127[22];
                    stage4_col127[27] <= stage3_col127[22];
                    stage4_col127[28] <= stage3_col127[22];
                    stage4_col127[29] <= stage3_col127[22];
                    stage4_col127[30] <= stage3_col127[22];
                    stage4_col127[31] <= stage3_col127[22];
                    stage4_col127[32] <= stage3_col127[22];
                    stage4_col127[33] <= stage3_col127[22];
                    stage4_col127[34] <= stage3_col127[22];
                    stage4_col127[35] <= stage3_col127[22];
                    stage4_col127[36] <= stage3_col127[22];
                    stage4_col127[37] <= stage3_col127[22];
                    stage4_col127[38] <= stage3_col127[22];
                    stage4_col127[39] <= stage3_col127[22];
                    stage4_col127[40] <= stage3_col127[22];
                    stage4_col127[41] <= stage3_col127[22];
                    stage4_col127[42] <= stage3_col127[22];
                    stage4_col127[43] <= stage3_col127[22];
                    stage4_col127[44] <= stage3_col127[22];
                    stage4_col127[45] <= stage3_col127[22];
                    stage4_col127[46] <= stage3_col127[22];
                    stage4_col127[47] <= stage3_col127[22];
                    stage4_col127[48] <= stage3_col127[22];
                    stage4_col127[49] <= stage3_col127[22];
                    stage4_col127[50] <= stage3_col127[22];
                    stage4_col127[51] <= stage3_col127[22];
                    stage4_col127[52] <= stage3_col127[22];
                    stage4_col127[53] <= stage3_col127[22];
                    stage4_col127[54] <= stage3_col127[22];
                    stage4_col127[55] <= stage3_col127[22];
                    stage4_col127[56] <= stage3_col127[22];
                end
            end
        end else begin : gen_stage4_no_pipe
            // Combinational assignment
            always_comb begin
                stage4_col0[0] = stage3_col0[0];
                stage4_col1[0] = stage3_col1[0];
                stage4_col2[0] = stage3_col2[0];
                stage4_col3[0] = ha_s3_c3_n0_s;
                stage4_col4[0] = ha_s3_c3_n0_c;
                stage4_col4[1] = stage3_col4[0];
                stage4_col5[0] = fa_s3_c5_n0_s;
                stage4_col6[0] = fa_s3_c5_n0_c;
                stage4_col6[1] = stage3_col6[0];
                stage4_col6[2] = stage3_col6[1];
                stage4_col7[0] = stage3_col7[0];
                stage4_col7[1] = stage3_col7[1];
                stage4_col8[0] = stage3_col8[0];
                stage4_col8[1] = stage3_col8[1];
                stage4_col9[0] = stage3_col9[0];
                stage4_col9[1] = stage3_col9[1];
                stage4_col10[0] = stage3_col10[0];
                stage4_col10[1] = stage3_col10[1];
                stage4_col11[0] = stage3_col11[0];
                stage4_col11[1] = stage3_col11[1];
                stage4_col12[0] = stage3_col12[0];
                stage4_col12[1] = stage3_col12[1];
                stage4_col13[0] = fa_s3_c13_n1_s;
                stage4_col13[1] = stage3_col13[3];
                stage4_col14[0] = fa_s3_c13_n1_c;
                stage4_col14[1] = fa_s3_c14_n2_s;
                stage4_col15[0] = fa_s3_c14_n2_c;
                stage4_col15[1] = fa_s3_c15_n3_s;
                stage4_col16[0] = fa_s3_c15_n3_c;
                stage4_col16[1] = fa_s3_c16_n4_s;
                stage4_col17[0] = fa_s3_c16_n4_c;
                stage4_col17[1] = fa_s3_c17_n5_s;
                stage4_col18[0] = fa_s3_c17_n5_c;
                stage4_col18[1] = fa_s3_c18_n6_s;
                stage4_col19[0] = fa_s3_c18_n6_c;
                stage4_col19[1] = fa_s3_c19_n7_s;
                stage4_col19[2] = stage3_col19[3];
                stage4_col19[3] = stage3_col19[4];
                stage4_col20[0] = fa_s3_c19_n7_c;
                stage4_col20[1] = fa_s3_c20_n8_s;
                stage4_col20[2] = stage3_col20[3];
                stage4_col21[0] = fa_s3_c20_n8_c;
                stage4_col21[1] = fa_s3_c21_n9_s;
                stage4_col21[2] = stage3_col21[3];
                stage4_col22[0] = fa_s3_c21_n9_c;
                stage4_col22[1] = fa_s3_c22_n10_s;
                stage4_col22[2] = stage3_col22[3];
                stage4_col23[0] = fa_s3_c22_n10_c;
                stage4_col23[1] = fa_s3_c23_n11_s;
                stage4_col23[2] = stage3_col23[3];
                stage4_col24[0] = fa_s3_c23_n11_c;
                stage4_col24[1] = fa_s3_c24_n12_s;
                stage4_col24[2] = stage3_col24[3];
                stage4_col25[0] = fa_s3_c24_n12_c;
                stage4_col25[1] = fa_s3_c25_n13_s;
                stage4_col25[2] = stage3_col25[3];
                stage4_col26[0] = fa_s3_c25_n13_c;
                stage4_col26[1] = fa_s3_c26_n14_s;
                stage4_col26[2] = stage3_col26[3];
                stage4_col27[0] = fa_s3_c26_n14_c;
                stage4_col27[1] = fa_s3_c27_n15_s;
                stage4_col27[2] = fa_s3_c27_n16_s;
                stage4_col28[0] = fa_s3_c27_n15_c;
                stage4_col28[1] = fa_s3_c27_n16_c;
                stage4_col28[2] = fa_s3_c28_n17_s;
                stage4_col28[3] = stage3_col28[3];
                stage4_col28[4] = stage3_col28[4];
                stage4_col29[0] = fa_s3_c28_n17_c;
                stage4_col29[1] = fa_s3_c29_n18_s;
                stage4_col29[2] = stage3_col29[3];
                stage4_col29[3] = stage3_col29[4];
                stage4_col30[0] = fa_s3_c29_n18_c;
                stage4_col30[1] = fa_s3_c30_n19_s;
                stage4_col30[2] = stage3_col30[3];
                stage4_col30[3] = stage3_col30[4];
                stage4_col31[0] = fa_s3_c30_n19_c;
                stage4_col31[1] = fa_s3_c31_n20_s;
                stage4_col31[2] = stage3_col31[3];
                stage4_col31[3] = stage3_col31[4];
                stage4_col32[0] = fa_s3_c31_n20_c;
                stage4_col32[1] = fa_s3_c32_n21_s;
                stage4_col32[2] = fa_s3_c32_n22_s;
                stage4_col32[3] = stage3_col32[6];
                stage4_col33[0] = fa_s3_c32_n21_c;
                stage4_col33[1] = fa_s3_c32_n22_c;
                stage4_col33[2] = fa_s3_c33_n23_s;
                stage4_col33[3] = fa_s3_c33_n24_s;
                stage4_col34[0] = fa_s3_c33_n23_c;
                stage4_col34[1] = fa_s3_c33_n24_c;
                stage4_col34[2] = fa_s3_c34_n25_s;
                stage4_col34[3] = fa_s3_c34_n26_s;
                stage4_col35[0] = fa_s3_c34_n25_c;
                stage4_col35[1] = fa_s3_c34_n26_c;
                stage4_col35[2] = fa_s3_c35_n27_s;
                stage4_col35[3] = fa_s3_c35_n28_s;
                stage4_col36[0] = fa_s3_c35_n27_c;
                stage4_col36[1] = fa_s3_c35_n28_c;
                stage4_col36[2] = fa_s3_c36_n29_s;
                stage4_col36[3] = fa_s3_c36_n30_s;
                stage4_col37[0] = fa_s3_c36_n29_c;
                stage4_col37[1] = fa_s3_c36_n30_c;
                stage4_col37[2] = fa_s3_c37_n31_s;
                stage4_col37[3] = fa_s3_c37_n32_s;
                stage4_col38[0] = fa_s3_c37_n31_c;
                stage4_col38[1] = fa_s3_c37_n32_c;
                stage4_col38[2] = fa_s3_c38_n33_s;
                stage4_col38[3] = fa_s3_c38_n34_s;
                stage4_col39[0] = fa_s3_c38_n33_c;
                stage4_col39[1] = fa_s3_c38_n34_c;
                stage4_col39[2] = fa_s3_c39_n35_s;
                stage4_col39[3] = fa_s3_c39_n36_s;
                stage4_col40[0] = fa_s3_c39_n35_c;
                stage4_col40[1] = fa_s3_c39_n36_c;
                stage4_col40[2] = fa_s3_c40_n37_s;
                stage4_col40[3] = fa_s3_c40_n38_s;
                stage4_col40[4] = stage3_col40[6];
                stage4_col40[5] = stage3_col40[7];
                stage4_col41[0] = fa_s3_c40_n37_c;
                stage4_col41[1] = fa_s3_c40_n38_c;
                stage4_col41[2] = fa_s3_c41_n39_s;
                stage4_col41[3] = fa_s3_c41_n40_s;
                stage4_col41[4] = stage3_col41[6];
                stage4_col42[0] = fa_s3_c41_n39_c;
                stage4_col42[1] = fa_s3_c41_n40_c;
                stage4_col42[2] = fa_s3_c42_n41_s;
                stage4_col42[3] = fa_s3_c42_n42_s;
                stage4_col42[4] = stage3_col42[6];
                stage4_col43[0] = fa_s3_c42_n41_c;
                stage4_col43[1] = fa_s3_c42_n42_c;
                stage4_col43[2] = fa_s3_c43_n43_s;
                stage4_col43[3] = fa_s3_c43_n44_s;
                stage4_col43[4] = stage3_col43[6];
                stage4_col44[0] = fa_s3_c43_n43_c;
                stage4_col44[1] = fa_s3_c43_n44_c;
                stage4_col44[2] = fa_s3_c44_n45_s;
                stage4_col44[3] = fa_s3_c44_n46_s;
                stage4_col44[4] = stage3_col44[6];
                stage4_col45[0] = fa_s3_c44_n45_c;
                stage4_col45[1] = fa_s3_c44_n46_c;
                stage4_col45[2] = fa_s3_c45_n47_s;
                stage4_col45[3] = fa_s3_c45_n48_s;
                stage4_col45[4] = stage3_col45[6];
                stage4_col46[0] = fa_s3_c45_n47_c;
                stage4_col46[1] = fa_s3_c45_n48_c;
                stage4_col46[2] = fa_s3_c46_n49_s;
                stage4_col46[3] = fa_s3_c46_n50_s;
                stage4_col46[4] = fa_s3_c46_n51_s;
                stage4_col47[0] = fa_s3_c46_n49_c;
                stage4_col47[1] = fa_s3_c46_n50_c;
                stage4_col47[2] = fa_s3_c46_n51_c;
                stage4_col47[3] = fa_s3_c47_n52_s;
                stage4_col47[4] = fa_s3_c47_n53_s;
                stage4_col47[5] = stage3_col47[6];
                stage4_col47[6] = stage3_col47[7];
                stage4_col48[0] = fa_s3_c47_n52_c;
                stage4_col48[1] = fa_s3_c47_n53_c;
                stage4_col48[2] = fa_s3_c48_n54_s;
                stage4_col48[3] = fa_s3_c48_n55_s;
                stage4_col48[4] = stage3_col48[6];
                stage4_col48[5] = stage3_col48[7];
                stage4_col49[0] = fa_s3_c48_n54_c;
                stage4_col49[1] = fa_s3_c48_n55_c;
                stage4_col49[2] = fa_s3_c49_n56_s;
                stage4_col49[3] = fa_s3_c49_n57_s;
                stage4_col49[4] = stage3_col49[6];
                stage4_col49[5] = stage3_col49[7];
                stage4_col50[0] = fa_s3_c49_n56_c;
                stage4_col50[1] = fa_s3_c49_n57_c;
                stage4_col50[2] = fa_s3_c50_n58_s;
                stage4_col50[3] = fa_s3_c50_n59_s;
                stage4_col50[4] = stage3_col50[6];
                stage4_col50[5] = stage3_col50[7];
                stage4_col51[0] = fa_s3_c50_n58_c;
                stage4_col51[1] = fa_s3_c50_n59_c;
                stage4_col51[2] = fa_s3_c51_n60_s;
                stage4_col51[3] = fa_s3_c51_n61_s;
                stage4_col51[4] = stage3_col51[6];
                stage4_col51[5] = stage3_col51[7];
                stage4_col52[0] = fa_s3_c51_n60_c;
                stage4_col52[1] = fa_s3_c51_n61_c;
                stage4_col52[2] = fa_s3_c52_n62_s;
                stage4_col52[3] = fa_s3_c52_n63_s;
                stage4_col52[4] = stage3_col52[6];
                stage4_col52[5] = stage3_col52[7];
                stage4_col53[0] = fa_s3_c52_n62_c;
                stage4_col53[1] = fa_s3_c52_n63_c;
                stage4_col53[2] = fa_s3_c53_n64_s;
                stage4_col53[3] = fa_s3_c53_n65_s;
                stage4_col53[4] = stage3_col53[6];
                stage4_col53[5] = stage3_col53[7];
                stage4_col54[0] = fa_s3_c53_n64_c;
                stage4_col54[1] = fa_s3_c53_n65_c;
                stage4_col54[2] = fa_s3_c54_n66_s;
                stage4_col54[3] = fa_s3_c54_n67_s;
                stage4_col54[4] = fa_s3_c54_n68_s;
                stage4_col54[5] = stage3_col54[9];
                stage4_col55[0] = fa_s3_c54_n66_c;
                stage4_col55[1] = fa_s3_c54_n67_c;
                stage4_col55[2] = fa_s3_c54_n68_c;
                stage4_col55[3] = fa_s3_c55_n69_s;
                stage4_col55[4] = fa_s3_c55_n70_s;
                stage4_col55[5] = fa_s3_c55_n71_s;
                stage4_col56[0] = fa_s3_c55_n69_c;
                stage4_col56[1] = fa_s3_c55_n70_c;
                stage4_col56[2] = fa_s3_c55_n71_c;
                stage4_col56[3] = fa_s3_c56_n72_s;
                stage4_col56[4] = fa_s3_c56_n73_s;
                stage4_col56[5] = fa_s3_c56_n74_s;
                stage4_col57[0] = fa_s3_c56_n72_c;
                stage4_col57[1] = fa_s3_c56_n73_c;
                stage4_col57[2] = fa_s3_c56_n74_c;
                stage4_col57[3] = fa_s3_c57_n75_s;
                stage4_col57[4] = fa_s3_c57_n76_s;
                stage4_col57[5] = fa_s3_c57_n77_s;
                stage4_col58[0] = fa_s3_c57_n75_c;
                stage4_col58[1] = fa_s3_c57_n76_c;
                stage4_col58[2] = fa_s3_c57_n77_c;
                stage4_col58[3] = fa_s3_c58_n78_s;
                stage4_col58[4] = fa_s3_c58_n79_s;
                stage4_col58[5] = fa_s3_c58_n80_s;
                stage4_col59[0] = fa_s3_c58_n78_c;
                stage4_col59[1] = fa_s3_c58_n79_c;
                stage4_col59[2] = fa_s3_c58_n80_c;
                stage4_col59[3] = fa_s3_c59_n81_s;
                stage4_col59[4] = fa_s3_c59_n82_s;
                stage4_col59[5] = fa_s3_c59_n83_s;
                stage4_col59[6] = stage3_col59[9];
                stage4_col59[7] = stage3_col59[10];
                stage4_col60[0] = fa_s3_c59_n81_c;
                stage4_col60[1] = fa_s3_c59_n82_c;
                stage4_col60[2] = fa_s3_c59_n83_c;
                stage4_col60[3] = fa_s3_c60_n84_s;
                stage4_col60[4] = fa_s3_c60_n85_s;
                stage4_col60[5] = fa_s3_c60_n86_s;
                stage4_col60[6] = stage3_col60[9];
                stage4_col61[0] = fa_s3_c60_n84_c;
                stage4_col61[1] = fa_s3_c60_n85_c;
                stage4_col61[2] = fa_s3_c60_n86_c;
                stage4_col61[3] = fa_s3_c61_n87_s;
                stage4_col61[4] = fa_s3_c61_n88_s;
                stage4_col61[5] = fa_s3_c61_n89_s;
                stage4_col61[6] = stage3_col61[9];
                stage4_col62[0] = fa_s3_c61_n87_c;
                stage4_col62[1] = fa_s3_c61_n88_c;
                stage4_col62[2] = fa_s3_c61_n89_c;
                stage4_col62[3] = fa_s3_c62_n90_s;
                stage4_col62[4] = fa_s3_c62_n91_s;
                stage4_col62[5] = fa_s3_c62_n92_s;
                stage4_col62[6] = stage3_col62[9];
                stage4_col63[0] = fa_s3_c62_n90_c;
                stage4_col63[1] = fa_s3_c62_n91_c;
                stage4_col63[2] = fa_s3_c62_n92_c;
                stage4_col63[3] = fa_s3_c63_n93_s;
                stage4_col63[4] = fa_s3_c63_n94_s;
                stage4_col63[5] = fa_s3_c63_n95_s;
                stage4_col63[6] = stage3_col63[9];
                stage4_col64[0] = fa_s3_c63_n93_c;
                stage4_col64[1] = fa_s3_c63_n94_c;
                stage4_col64[2] = fa_s3_c63_n95_c;
                stage4_col64[3] = fa_s3_c64_n96_s;
                stage4_col64[4] = fa_s3_c64_n97_s;
                stage4_col64[5] = fa_s3_c64_n98_s;
                stage4_col64[6] = stage3_col64[9];
                stage4_col64[7] = stage3_col64[10];
                stage4_col65[0] = fa_s3_c64_n96_c;
                stage4_col65[1] = fa_s3_c64_n97_c;
                stage4_col65[2] = fa_s3_c64_n98_c;
                stage4_col65[3] = fa_s3_c65_n99_s;
                stage4_col65[4] = fa_s3_c65_n100_s;
                stage4_col65[5] = fa_s3_c65_n101_s;
                stage4_col65[6] = stage3_col65[9];
                stage4_col66[0] = fa_s3_c65_n99_c;
                stage4_col66[1] = fa_s3_c65_n100_c;
                stage4_col66[2] = fa_s3_c65_n101_c;
                stage4_col66[3] = fa_s3_c66_n102_s;
                stage4_col66[4] = fa_s3_c66_n103_s;
                stage4_col66[5] = fa_s3_c66_n104_s;
                stage4_col66[6] = stage3_col66[9];
                stage4_col66[7] = stage3_col66[10];
                stage4_col67[0] = fa_s3_c66_n102_c;
                stage4_col67[1] = fa_s3_c66_n103_c;
                stage4_col67[2] = fa_s3_c66_n104_c;
                stage4_col67[3] = fa_s3_c67_n105_s;
                stage4_col67[4] = fa_s3_c67_n106_s;
                stage4_col67[5] = fa_s3_c67_n107_s;
                stage4_col67[6] = stage3_col67[9];
                stage4_col68[0] = fa_s3_c67_n105_c;
                stage4_col68[1] = fa_s3_c67_n106_c;
                stage4_col68[2] = fa_s3_c67_n107_c;
                stage4_col68[3] = fa_s3_c68_n108_s;
                stage4_col68[4] = fa_s3_c68_n109_s;
                stage4_col68[5] = fa_s3_c68_n110_s;
                stage4_col68[6] = stage3_col68[9];
                stage4_col68[7] = stage3_col68[10];
                stage4_col69[0] = fa_s3_c68_n108_c;
                stage4_col69[1] = fa_s3_c68_n109_c;
                stage4_col69[2] = fa_s3_c68_n110_c;
                stage4_col69[3] = fa_s3_c69_n111_s;
                stage4_col69[4] = fa_s3_c69_n112_s;
                stage4_col69[5] = fa_s3_c69_n113_s;
                stage4_col69[6] = stage3_col69[9];
                stage4_col70[0] = fa_s3_c69_n111_c;
                stage4_col70[1] = fa_s3_c69_n112_c;
                stage4_col70[2] = fa_s3_c69_n113_c;
                stage4_col70[3] = fa_s3_c70_n114_s;
                stage4_col70[4] = fa_s3_c70_n115_s;
                stage4_col70[5] = fa_s3_c70_n116_s;
                stage4_col70[6] = stage3_col70[9];
                stage4_col70[7] = stage3_col70[10];
                stage4_col71[0] = fa_s3_c70_n114_c;
                stage4_col71[1] = fa_s3_c70_n115_c;
                stage4_col71[2] = fa_s3_c70_n116_c;
                stage4_col71[3] = fa_s3_c71_n117_s;
                stage4_col71[4] = fa_s3_c71_n118_s;
                stage4_col71[5] = fa_s3_c71_n119_s;
                stage4_col71[6] = stage3_col71[9];
                stage4_col72[0] = fa_s3_c71_n117_c;
                stage4_col72[1] = fa_s3_c71_n118_c;
                stage4_col72[2] = fa_s3_c71_n119_c;
                stage4_col72[3] = fa_s3_c72_n120_s;
                stage4_col72[4] = fa_s3_c72_n121_s;
                stage4_col72[5] = fa_s3_c72_n122_s;
                stage4_col72[6] = stage3_col72[9];
                stage4_col72[7] = stage3_col72[10];
                stage4_col73[0] = fa_s3_c72_n120_c;
                stage4_col73[1] = fa_s3_c72_n121_c;
                stage4_col73[2] = fa_s3_c72_n122_c;
                stage4_col73[3] = fa_s3_c73_n123_s;
                stage4_col73[4] = fa_s3_c73_n124_s;
                stage4_col73[5] = fa_s3_c73_n125_s;
                stage4_col73[6] = stage3_col73[9];
                stage4_col74[0] = fa_s3_c73_n123_c;
                stage4_col74[1] = fa_s3_c73_n124_c;
                stage4_col74[2] = fa_s3_c73_n125_c;
                stage4_col74[3] = fa_s3_c74_n126_s;
                stage4_col74[4] = fa_s3_c74_n127_s;
                stage4_col74[5] = fa_s3_c74_n128_s;
                stage4_col74[6] = stage3_col74[9];
                stage4_col74[7] = stage3_col74[10];
                stage4_col75[0] = fa_s3_c74_n126_c;
                stage4_col75[1] = fa_s3_c74_n127_c;
                stage4_col75[2] = fa_s3_c74_n128_c;
                stage4_col75[3] = fa_s3_c75_n129_s;
                stage4_col75[4] = fa_s3_c75_n130_s;
                stage4_col75[5] = fa_s3_c75_n131_s;
                stage4_col75[6] = stage3_col75[9];
                stage4_col76[0] = fa_s3_c75_n129_c;
                stage4_col76[1] = fa_s3_c75_n130_c;
                stage4_col76[2] = fa_s3_c75_n131_c;
                stage4_col76[3] = fa_s3_c76_n132_s;
                stage4_col76[4] = fa_s3_c76_n133_s;
                stage4_col76[5] = fa_s3_c76_n134_s;
                stage4_col76[6] = stage3_col76[9];
                stage4_col76[7] = stage3_col76[10];
                stage4_col77[0] = fa_s3_c76_n132_c;
                stage4_col77[1] = fa_s3_c76_n133_c;
                stage4_col77[2] = fa_s3_c76_n134_c;
                stage4_col77[3] = fa_s3_c77_n135_s;
                stage4_col77[4] = fa_s3_c77_n136_s;
                stage4_col77[5] = fa_s3_c77_n137_s;
                stage4_col77[6] = stage3_col77[9];
                stage4_col78[0] = fa_s3_c77_n135_c;
                stage4_col78[1] = fa_s3_c77_n136_c;
                stage4_col78[2] = fa_s3_c77_n137_c;
                stage4_col78[3] = fa_s3_c78_n138_s;
                stage4_col78[4] = fa_s3_c78_n139_s;
                stage4_col78[5] = fa_s3_c78_n140_s;
                stage4_col78[6] = stage3_col78[9];
                stage4_col78[7] = stage3_col78[10];
                stage4_col79[0] = fa_s3_c78_n138_c;
                stage4_col79[1] = fa_s3_c78_n139_c;
                stage4_col79[2] = fa_s3_c78_n140_c;
                stage4_col79[3] = fa_s3_c79_n141_s;
                stage4_col79[4] = fa_s3_c79_n142_s;
                stage4_col79[5] = fa_s3_c79_n143_s;
                stage4_col79[6] = stage3_col79[9];
                stage4_col80[0] = fa_s3_c79_n141_c;
                stage4_col80[1] = fa_s3_c79_n142_c;
                stage4_col80[2] = fa_s3_c79_n143_c;
                stage4_col80[3] = fa_s3_c80_n144_s;
                stage4_col80[4] = fa_s3_c80_n145_s;
                stage4_col80[5] = fa_s3_c80_n146_s;
                stage4_col80[6] = stage3_col80[9];
                stage4_col80[7] = stage3_col80[10];
                stage4_col81[0] = fa_s3_c80_n144_c;
                stage4_col81[1] = fa_s3_c80_n145_c;
                stage4_col81[2] = fa_s3_c80_n146_c;
                stage4_col81[3] = fa_s3_c81_n147_s;
                stage4_col81[4] = fa_s3_c81_n148_s;
                stage4_col81[5] = fa_s3_c81_n149_s;
                stage4_col81[6] = stage3_col81[9];
                stage4_col82[0] = fa_s3_c81_n147_c;
                stage4_col82[1] = fa_s3_c81_n148_c;
                stage4_col82[2] = fa_s3_c81_n149_c;
                stage4_col82[3] = fa_s3_c82_n150_s;
                stage4_col82[4] = fa_s3_c82_n151_s;
                stage4_col82[5] = fa_s3_c82_n152_s;
                stage4_col82[6] = stage3_col82[9];
                stage4_col82[7] = stage3_col82[10];
                stage4_col83[0] = fa_s3_c82_n150_c;
                stage4_col83[1] = fa_s3_c82_n151_c;
                stage4_col83[2] = fa_s3_c82_n152_c;
                stage4_col83[3] = fa_s3_c83_n153_s;
                stage4_col83[4] = fa_s3_c83_n154_s;
                stage4_col83[5] = fa_s3_c83_n155_s;
                stage4_col83[6] = stage3_col83[9];
                stage4_col84[0] = fa_s3_c83_n153_c;
                stage4_col84[1] = fa_s3_c83_n154_c;
                stage4_col84[2] = fa_s3_c83_n155_c;
                stage4_col84[3] = fa_s3_c84_n156_s;
                stage4_col84[4] = fa_s3_c84_n157_s;
                stage4_col84[5] = fa_s3_c84_n158_s;
                stage4_col84[6] = stage3_col84[9];
                stage4_col84[7] = stage3_col84[10];
                stage4_col85[0] = fa_s3_c84_n156_c;
                stage4_col85[1] = fa_s3_c84_n157_c;
                stage4_col85[2] = fa_s3_c84_n158_c;
                stage4_col85[3] = fa_s3_c85_n159_s;
                stage4_col85[4] = fa_s3_c85_n160_s;
                stage4_col85[5] = fa_s3_c85_n161_s;
                stage4_col85[6] = stage3_col85[9];
                stage4_col86[0] = fa_s3_c85_n159_c;
                stage4_col86[1] = fa_s3_c85_n160_c;
                stage4_col86[2] = fa_s3_c85_n161_c;
                stage4_col86[3] = fa_s3_c86_n162_s;
                stage4_col86[4] = fa_s3_c86_n163_s;
                stage4_col86[5] = fa_s3_c86_n164_s;
                stage4_col86[6] = stage3_col86[9];
                stage4_col86[7] = stage3_col86[10];
                stage4_col87[0] = fa_s3_c86_n162_c;
                stage4_col87[1] = fa_s3_c86_n163_c;
                stage4_col87[2] = fa_s3_c86_n164_c;
                stage4_col87[3] = fa_s3_c87_n165_s;
                stage4_col87[4] = fa_s3_c87_n166_s;
                stage4_col87[5] = fa_s3_c87_n167_s;
                stage4_col87[6] = stage3_col87[9];
                stage4_col88[0] = fa_s3_c87_n165_c;
                stage4_col88[1] = fa_s3_c87_n166_c;
                stage4_col88[2] = fa_s3_c87_n167_c;
                stage4_col88[3] = fa_s3_c88_n168_s;
                stage4_col88[4] = fa_s3_c88_n169_s;
                stage4_col88[5] = fa_s3_c88_n170_s;
                stage4_col88[6] = stage3_col88[9];
                stage4_col88[7] = stage3_col88[10];
                stage4_col89[0] = fa_s3_c88_n168_c;
                stage4_col89[1] = fa_s3_c88_n169_c;
                stage4_col89[2] = fa_s3_c88_n170_c;
                stage4_col89[3] = fa_s3_c89_n171_s;
                stage4_col89[4] = fa_s3_c89_n172_s;
                stage4_col89[5] = fa_s3_c89_n173_s;
                stage4_col89[6] = stage3_col89[9];
                stage4_col90[0] = fa_s3_c89_n171_c;
                stage4_col90[1] = fa_s3_c89_n172_c;
                stage4_col90[2] = fa_s3_c89_n173_c;
                stage4_col90[3] = fa_s3_c90_n174_s;
                stage4_col90[4] = fa_s3_c90_n175_s;
                stage4_col90[5] = fa_s3_c90_n176_s;
                stage4_col90[6] = stage3_col90[9];
                stage4_col90[7] = stage3_col90[10];
                stage4_col91[0] = fa_s3_c90_n174_c;
                stage4_col91[1] = fa_s3_c90_n175_c;
                stage4_col91[2] = fa_s3_c90_n176_c;
                stage4_col91[3] = fa_s3_c91_n177_s;
                stage4_col91[4] = fa_s3_c91_n178_s;
                stage4_col91[5] = fa_s3_c91_n179_s;
                stage4_col91[6] = stage3_col91[9];
                stage4_col92[0] = fa_s3_c91_n177_c;
                stage4_col92[1] = fa_s3_c91_n178_c;
                stage4_col92[2] = fa_s3_c91_n179_c;
                stage4_col92[3] = fa_s3_c92_n180_s;
                stage4_col92[4] = fa_s3_c92_n181_s;
                stage4_col92[5] = fa_s3_c92_n182_s;
                stage4_col92[6] = stage3_col92[9];
                stage4_col92[7] = stage3_col92[10];
                stage4_col93[0] = fa_s3_c92_n180_c;
                stage4_col93[1] = fa_s3_c92_n181_c;
                stage4_col93[2] = fa_s3_c92_n182_c;
                stage4_col93[3] = fa_s3_c93_n183_s;
                stage4_col93[4] = fa_s3_c93_n184_s;
                stage4_col93[5] = fa_s3_c93_n185_s;
                stage4_col93[6] = stage3_col93[9];
                stage4_col94[0] = fa_s3_c93_n183_c;
                stage4_col94[1] = fa_s3_c93_n184_c;
                stage4_col94[2] = fa_s3_c93_n185_c;
                stage4_col94[3] = fa_s3_c94_n186_s;
                stage4_col94[4] = fa_s3_c94_n187_s;
                stage4_col94[5] = fa_s3_c94_n188_s;
                stage4_col94[6] = stage3_col94[9];
                stage4_col94[7] = stage3_col94[10];
                stage4_col95[0] = fa_s3_c94_n186_c;
                stage4_col95[1] = fa_s3_c94_n187_c;
                stage4_col95[2] = fa_s3_c94_n188_c;
                stage4_col95[3] = fa_s3_c95_n189_s;
                stage4_col95[4] = fa_s3_c95_n190_s;
                stage4_col95[5] = fa_s3_c95_n191_s;
                stage4_col95[6] = stage3_col95[9];
                stage4_col96[0] = fa_s3_c95_n189_c;
                stage4_col96[1] = fa_s3_c95_n190_c;
                stage4_col96[2] = fa_s3_c95_n191_c;
                stage4_col96[3] = fa_s3_c96_n192_s;
                stage4_col96[4] = fa_s3_c96_n193_s;
                stage4_col96[5] = fa_s3_c96_n194_s;
                stage4_col96[6] = stage3_col96[9];
                stage4_col96[7] = stage3_col96[10];
                stage4_col97[0] = fa_s3_c96_n192_c;
                stage4_col97[1] = fa_s3_c96_n193_c;
                stage4_col97[2] = fa_s3_c96_n194_c;
                stage4_col97[3] = fa_s3_c97_n195_s;
                stage4_col97[4] = fa_s3_c97_n196_s;
                stage4_col97[5] = fa_s3_c97_n197_s;
                stage4_col97[6] = stage3_col97[9];
                stage4_col98[0] = fa_s3_c97_n195_c;
                stage4_col98[1] = fa_s3_c97_n196_c;
                stage4_col98[2] = fa_s3_c97_n197_c;
                stage4_col98[3] = fa_s3_c98_n198_s;
                stage4_col98[4] = fa_s3_c98_n199_s;
                stage4_col98[5] = fa_s3_c98_n200_s;
                stage4_col98[6] = stage3_col98[9];
                stage4_col98[7] = stage3_col98[10];
                stage4_col99[0] = fa_s3_c98_n198_c;
                stage4_col99[1] = fa_s3_c98_n199_c;
                stage4_col99[2] = fa_s3_c98_n200_c;
                stage4_col99[3] = fa_s3_c99_n201_s;
                stage4_col99[4] = fa_s3_c99_n202_s;
                stage4_col99[5] = fa_s3_c99_n203_s;
                stage4_col99[6] = stage3_col99[9];
                stage4_col100[0] = fa_s3_c99_n201_c;
                stage4_col100[1] = fa_s3_c99_n202_c;
                stage4_col100[2] = fa_s3_c99_n203_c;
                stage4_col100[3] = fa_s3_c100_n204_s;
                stage4_col100[4] = fa_s3_c100_n205_s;
                stage4_col100[5] = fa_s3_c100_n206_s;
                stage4_col100[6] = stage3_col100[9];
                stage4_col100[7] = stage3_col100[10];
                stage4_col101[0] = fa_s3_c100_n204_c;
                stage4_col101[1] = fa_s3_c100_n205_c;
                stage4_col101[2] = fa_s3_c100_n206_c;
                stage4_col101[3] = fa_s3_c101_n207_s;
                stage4_col101[4] = fa_s3_c101_n208_s;
                stage4_col101[5] = fa_s3_c101_n209_s;
                stage4_col101[6] = stage3_col101[9];
                stage4_col102[0] = fa_s3_c101_n207_c;
                stage4_col102[1] = fa_s3_c101_n208_c;
                stage4_col102[2] = fa_s3_c101_n209_c;
                stage4_col102[3] = fa_s3_c102_n210_s;
                stage4_col102[4] = fa_s3_c102_n211_s;
                stage4_col102[5] = fa_s3_c102_n212_s;
                stage4_col102[6] = stage3_col102[9];
                stage4_col102[7] = stage3_col102[10];
                stage4_col103[0] = fa_s3_c102_n210_c;
                stage4_col103[1] = fa_s3_c102_n211_c;
                stage4_col103[2] = fa_s3_c102_n212_c;
                stage4_col103[3] = fa_s3_c103_n213_s;
                stage4_col103[4] = fa_s3_c103_n214_s;
                stage4_col103[5] = fa_s3_c103_n215_s;
                stage4_col103[6] = stage3_col103[9];
                stage4_col104[0] = fa_s3_c103_n213_c;
                stage4_col104[1] = fa_s3_c103_n214_c;
                stage4_col104[2] = fa_s3_c103_n215_c;
                stage4_col104[3] = fa_s3_c104_n216_s;
                stage4_col104[4] = fa_s3_c104_n217_s;
                stage4_col104[5] = fa_s3_c104_n218_s;
                stage4_col104[6] = stage3_col104[9];
                stage4_col104[7] = stage3_col104[10];
                stage4_col105[0] = fa_s3_c104_n216_c;
                stage4_col105[1] = fa_s3_c104_n217_c;
                stage4_col105[2] = fa_s3_c104_n218_c;
                stage4_col105[3] = fa_s3_c105_n219_s;
                stage4_col105[4] = fa_s3_c105_n220_s;
                stage4_col105[5] = fa_s3_c105_n221_s;
                stage4_col105[6] = stage3_col105[9];
                stage4_col106[0] = fa_s3_c105_n219_c;
                stage4_col106[1] = fa_s3_c105_n220_c;
                stage4_col106[2] = fa_s3_c105_n221_c;
                stage4_col106[3] = fa_s3_c106_n222_s;
                stage4_col106[4] = fa_s3_c106_n223_s;
                stage4_col106[5] = fa_s3_c106_n224_s;
                stage4_col106[6] = stage3_col106[9];
                stage4_col106[7] = stage3_col106[10];
                stage4_col107[0] = fa_s3_c106_n222_c;
                stage4_col107[1] = fa_s3_c106_n223_c;
                stage4_col107[2] = fa_s3_c106_n224_c;
                stage4_col107[3] = fa_s3_c107_n225_s;
                stage4_col107[4] = fa_s3_c107_n226_s;
                stage4_col107[5] = fa_s3_c107_n227_s;
                stage4_col107[6] = stage3_col107[9];
                stage4_col108[0] = fa_s3_c107_n225_c;
                stage4_col108[1] = fa_s3_c107_n226_c;
                stage4_col108[2] = fa_s3_c107_n227_c;
                stage4_col108[3] = fa_s3_c108_n228_s;
                stage4_col108[4] = fa_s3_c108_n229_s;
                stage4_col108[5] = fa_s3_c108_n230_s;
                stage4_col108[6] = stage3_col108[9];
                stage4_col108[7] = stage3_col108[10];
                stage4_col109[0] = fa_s3_c108_n228_c;
                stage4_col109[1] = fa_s3_c108_n229_c;
                stage4_col109[2] = fa_s3_c108_n230_c;
                stage4_col109[3] = fa_s3_c109_n231_s;
                stage4_col109[4] = fa_s3_c109_n232_s;
                stage4_col109[5] = fa_s3_c109_n233_s;
                stage4_col109[6] = stage3_col109[9];
                stage4_col110[0] = fa_s3_c109_n231_c;
                stage4_col110[1] = fa_s3_c109_n232_c;
                stage4_col110[2] = fa_s3_c109_n233_c;
                stage4_col110[3] = fa_s3_c110_n234_s;
                stage4_col110[4] = fa_s3_c110_n235_s;
                stage4_col110[5] = fa_s3_c110_n236_s;
                stage4_col110[6] = stage3_col110[9];
                stage4_col110[7] = stage3_col110[10];
                stage4_col111[0] = fa_s3_c110_n234_c;
                stage4_col111[1] = fa_s3_c110_n235_c;
                stage4_col111[2] = fa_s3_c110_n236_c;
                stage4_col111[3] = fa_s3_c111_n237_s;
                stage4_col111[4] = fa_s3_c111_n238_s;
                stage4_col111[5] = fa_s3_c111_n239_s;
                stage4_col111[6] = stage3_col111[9];
                stage4_col112[0] = fa_s3_c111_n237_c;
                stage4_col112[1] = fa_s3_c111_n238_c;
                stage4_col112[2] = fa_s3_c111_n239_c;
                stage4_col112[3] = fa_s3_c112_n240_s;
                stage4_col112[4] = fa_s3_c112_n241_s;
                stage4_col112[5] = fa_s3_c112_n242_s;
                stage4_col112[6] = stage3_col112[9];
                stage4_col112[7] = stage3_col112[10];
                stage4_col113[0] = fa_s3_c112_n240_c;
                stage4_col113[1] = fa_s3_c112_n241_c;
                stage4_col113[2] = fa_s3_c112_n242_c;
                stage4_col113[3] = fa_s3_c113_n243_s;
                stage4_col113[4] = fa_s3_c113_n244_s;
                stage4_col113[5] = fa_s3_c113_n245_s;
                stage4_col113[6] = stage3_col113[9];
                stage4_col114[0] = fa_s3_c113_n243_c;
                stage4_col114[1] = fa_s3_c113_n244_c;
                stage4_col114[2] = fa_s3_c113_n245_c;
                stage4_col114[3] = fa_s3_c114_n246_s;
                stage4_col114[4] = fa_s3_c114_n247_s;
                stage4_col114[5] = fa_s3_c114_n248_s;
                stage4_col114[6] = stage3_col114[9];
                stage4_col114[7] = stage3_col114[10];
                stage4_col115[0] = fa_s3_c114_n246_c;
                stage4_col115[1] = fa_s3_c114_n247_c;
                stage4_col115[2] = fa_s3_c114_n248_c;
                stage4_col115[3] = fa_s3_c115_n249_s;
                stage4_col115[4] = fa_s3_c115_n250_s;
                stage4_col115[5] = fa_s3_c115_n251_s;
                stage4_col115[6] = stage3_col115[9];
                stage4_col116[0] = fa_s3_c115_n249_c;
                stage4_col116[1] = fa_s3_c115_n250_c;
                stage4_col116[2] = fa_s3_c115_n251_c;
                stage4_col116[3] = fa_s3_c116_n252_s;
                stage4_col116[4] = fa_s3_c116_n253_s;
                stage4_col116[5] = fa_s3_c116_n254_s;
                stage4_col116[6] = stage3_col116[9];
                stage4_col116[7] = stage3_col116[10];
                stage4_col117[0] = fa_s3_c116_n252_c;
                stage4_col117[1] = fa_s3_c116_n253_c;
                stage4_col117[2] = fa_s3_c116_n254_c;
                stage4_col117[3] = fa_s3_c117_n255_s;
                stage4_col117[4] = fa_s3_c117_n256_s;
                stage4_col117[5] = fa_s3_c117_n257_s;
                stage4_col117[6] = stage3_col117[9];
                stage4_col118[0] = fa_s3_c117_n255_c;
                stage4_col118[1] = fa_s3_c117_n256_c;
                stage4_col118[2] = fa_s3_c117_n257_c;
                stage4_col118[3] = fa_s3_c118_n258_s;
                stage4_col118[4] = fa_s3_c118_n259_s;
                stage4_col118[5] = fa_s3_c118_n260_s;
                stage4_col118[6] = stage3_col118[9];
                stage4_col118[7] = stage3_col118[10];
                stage4_col119[0] = fa_s3_c118_n258_c;
                stage4_col119[1] = fa_s3_c118_n259_c;
                stage4_col119[2] = fa_s3_c118_n260_c;
                stage4_col119[3] = fa_s3_c119_n261_s;
                stage4_col119[4] = fa_s3_c119_n262_s;
                stage4_col119[5] = fa_s3_c119_n263_s;
                stage4_col119[6] = stage3_col119[9];
                stage4_col120[0] = fa_s3_c119_n261_c;
                stage4_col120[1] = fa_s3_c119_n262_c;
                stage4_col120[2] = fa_s3_c119_n263_c;
                stage4_col120[3] = fa_s3_c120_n264_s;
                stage4_col120[4] = fa_s3_c120_n265_s;
                stage4_col120[5] = fa_s3_c120_n266_s;
                stage4_col120[6] = stage3_col120[9];
                stage4_col120[7] = stage3_col120[10];
                stage4_col121[0] = fa_s3_c120_n264_c;
                stage4_col121[1] = fa_s3_c120_n265_c;
                stage4_col121[2] = fa_s3_c120_n266_c;
                stage4_col121[3] = fa_s3_c121_n267_s;
                stage4_col121[4] = fa_s3_c121_n268_s;
                stage4_col121[5] = fa_s3_c121_n269_s;
                stage4_col121[6] = stage3_col121[9];
                stage4_col122[0] = fa_s3_c121_n267_c;
                stage4_col122[1] = fa_s3_c121_n268_c;
                stage4_col122[2] = fa_s3_c121_n269_c;
                stage4_col122[3] = fa_s3_c122_n270_s;
                stage4_col122[4] = fa_s3_c122_n271_s;
                stage4_col122[5] = fa_s3_c122_n272_s;
                stage4_col122[6] = stage3_col122[9];
                stage4_col122[7] = stage3_col122[10];
                stage4_col123[0] = fa_s3_c122_n270_c;
                stage4_col123[1] = fa_s3_c122_n271_c;
                stage4_col123[2] = fa_s3_c122_n272_c;
                stage4_col123[3] = fa_s3_c123_n273_s;
                stage4_col123[4] = fa_s3_c123_n274_s;
                stage4_col123[5] = fa_s3_c123_n275_s;
                stage4_col123[6] = stage3_col123[9];
                stage4_col124[0] = fa_s3_c123_n273_c;
                stage4_col124[1] = fa_s3_c123_n274_c;
                stage4_col124[2] = fa_s3_c123_n275_c;
                stage4_col124[3] = fa_s3_c124_n276_s;
                stage4_col124[4] = fa_s3_c124_n277_s;
                stage4_col124[5] = fa_s3_c124_n278_s;
                stage4_col124[6] = stage3_col124[9];
                stage4_col124[7] = stage3_col124[10];
                stage4_col125[0] = fa_s3_c124_n276_c;
                stage4_col125[1] = fa_s3_c124_n277_c;
                stage4_col125[2] = fa_s3_c124_n278_c;
                stage4_col125[3] = fa_s3_c125_n279_s;
                stage4_col125[4] = fa_s3_c125_n280_s;
                stage4_col125[5] = fa_s3_c125_n281_s;
                stage4_col125[6] = stage3_col125[9];
                stage4_col126[0] = fa_s3_c125_n279_c;
                stage4_col126[1] = fa_s3_c125_n280_c;
                stage4_col126[2] = fa_s3_c125_n281_c;
                stage4_col126[3] = fa_s3_c126_n282_s;
                stage4_col126[4] = fa_s3_c126_n283_s;
                stage4_col126[5] = fa_s3_c126_n284_s;
                stage4_col126[6] = stage3_col126[9];
                stage4_col126[7] = stage3_col126[10];
                stage4_col127[0] = fa_s3_c126_n282_c;
                stage4_col127[1] = fa_s3_c126_n283_c;
                stage4_col127[2] = fa_s3_c126_n284_c;
                stage4_col127[3] = stage3_col127[0];
                stage4_col127[4] = stage3_col127[1];
                stage4_col127[5] = stage3_col127[2];
                stage4_col127[6] = stage3_col127[3];
                stage4_col127[7] = stage3_col127[4];
                stage4_col127[8] = stage3_col127[5];
                stage4_col127[9] = stage3_col127[6];
                stage4_col127[10] = stage3_col127[7];
                stage4_col127[11] = stage3_col127[8];
                stage4_col127[12] = stage3_col127[9];
                stage4_col127[13] = stage3_col127[10];
                stage4_col127[14] = stage3_col127[11];
                stage4_col127[15] = stage3_col127[12];
                stage4_col127[16] = stage3_col127[13];
                stage4_col127[17] = stage3_col127[14];
                stage4_col127[18] = stage3_col127[15];
                stage4_col127[19] = stage3_col127[16];
                stage4_col127[20] = stage3_col127[17];
                stage4_col127[21] = stage3_col127[18];
                stage4_col127[22] = stage3_col127[19];
                stage4_col127[23] = stage3_col127[20];
                stage4_col127[24] = stage3_col127[21];
                stage4_col127[25] = stage3_col127[22];
                stage4_col127[26] = stage3_col127[22];
                stage4_col127[27] = stage3_col127[22];
                stage4_col127[28] = stage3_col127[22];
                stage4_col127[29] = stage3_col127[22];
                stage4_col127[30] = stage3_col127[22];
                stage4_col127[31] = stage3_col127[22];
                stage4_col127[32] = stage3_col127[22];
                stage4_col127[33] = stage3_col127[22];
                stage4_col127[34] = stage3_col127[22];
                stage4_col127[35] = stage3_col127[22];
                stage4_col127[36] = stage3_col127[22];
                stage4_col127[37] = stage3_col127[22];
                stage4_col127[38] = stage3_col127[22];
                stage4_col127[39] = stage3_col127[22];
                stage4_col127[40] = stage3_col127[22];
                stage4_col127[41] = stage3_col127[22];
                stage4_col127[42] = stage3_col127[22];
                stage4_col127[43] = stage3_col127[22];
                stage4_col127[44] = stage3_col127[22];
                stage4_col127[45] = stage3_col127[22];
                stage4_col127[46] = stage3_col127[22];
                stage4_col127[47] = stage3_col127[22];
                stage4_col127[48] = stage3_col127[22];
                stage4_col127[49] = stage3_col127[22];
                stage4_col127[50] = stage3_col127[22];
                stage4_col127[51] = stage3_col127[22];
                stage4_col127[52] = stage3_col127[22];
                stage4_col127[53] = stage3_col127[22];
                stage4_col127[54] = stage3_col127[22];
                stage4_col127[55] = stage3_col127[22];
                stage4_col127[56] = stage3_col127[22];
            end
        end
    endgenerate

    // Stage 5: Reduction
    fa fa_s4_c6_n0 (
        .a(stage4_col6[0]),
        .b(stage4_col6[1]),
        .c_in(stage4_col6[2]),
        .s(fa_s4_c6_n0_s),
        .c_out(fa_s4_c6_n0_c)
    );

    fa fa_s4_c19_n1 (
        .a(stage4_col19[0]),
        .b(stage4_col19[1]),
        .c_in(stage4_col19[2]),
        .s(fa_s4_c19_n1_s),
        .c_out(fa_s4_c19_n1_c)
    );

    fa fa_s4_c20_n2 (
        .a(stage4_col20[0]),
        .b(stage4_col20[1]),
        .c_in(stage4_col20[2]),
        .s(fa_s4_c20_n2_s),
        .c_out(fa_s4_c20_n2_c)
    );

    fa fa_s4_c21_n3 (
        .a(stage4_col21[0]),
        .b(stage4_col21[1]),
        .c_in(stage4_col21[2]),
        .s(fa_s4_c21_n3_s),
        .c_out(fa_s4_c21_n3_c)
    );

    fa fa_s4_c22_n4 (
        .a(stage4_col22[0]),
        .b(stage4_col22[1]),
        .c_in(stage4_col22[2]),
        .s(fa_s4_c22_n4_s),
        .c_out(fa_s4_c22_n4_c)
    );

    fa fa_s4_c23_n5 (
        .a(stage4_col23[0]),
        .b(stage4_col23[1]),
        .c_in(stage4_col23[2]),
        .s(fa_s4_c23_n5_s),
        .c_out(fa_s4_c23_n5_c)
    );

    fa fa_s4_c24_n6 (
        .a(stage4_col24[0]),
        .b(stage4_col24[1]),
        .c_in(stage4_col24[2]),
        .s(fa_s4_c24_n6_s),
        .c_out(fa_s4_c24_n6_c)
    );

    fa fa_s4_c25_n7 (
        .a(stage4_col25[0]),
        .b(stage4_col25[1]),
        .c_in(stage4_col25[2]),
        .s(fa_s4_c25_n7_s),
        .c_out(fa_s4_c25_n7_c)
    );

    fa fa_s4_c26_n8 (
        .a(stage4_col26[0]),
        .b(stage4_col26[1]),
        .c_in(stage4_col26[2]),
        .s(fa_s4_c26_n8_s),
        .c_out(fa_s4_c26_n8_c)
    );

    fa fa_s4_c27_n9 (
        .a(stage4_col27[0]),
        .b(stage4_col27[1]),
        .c_in(stage4_col27[2]),
        .s(fa_s4_c27_n9_s),
        .c_out(fa_s4_c27_n9_c)
    );

    fa fa_s4_c28_n10 (
        .a(stage4_col28[0]),
        .b(stage4_col28[1]),
        .c_in(stage4_col28[2]),
        .s(fa_s4_c28_n10_s),
        .c_out(fa_s4_c28_n10_c)
    );

    fa fa_s4_c29_n11 (
        .a(stage4_col29[0]),
        .b(stage4_col29[1]),
        .c_in(stage4_col29[2]),
        .s(fa_s4_c29_n11_s),
        .c_out(fa_s4_c29_n11_c)
    );

    fa fa_s4_c30_n12 (
        .a(stage4_col30[0]),
        .b(stage4_col30[1]),
        .c_in(stage4_col30[2]),
        .s(fa_s4_c30_n12_s),
        .c_out(fa_s4_c30_n12_c)
    );

    fa fa_s4_c31_n13 (
        .a(stage4_col31[0]),
        .b(stage4_col31[1]),
        .c_in(stage4_col31[2]),
        .s(fa_s4_c31_n13_s),
        .c_out(fa_s4_c31_n13_c)
    );

    fa fa_s4_c32_n14 (
        .a(stage4_col32[0]),
        .b(stage4_col32[1]),
        .c_in(stage4_col32[2]),
        .s(fa_s4_c32_n14_s),
        .c_out(fa_s4_c32_n14_c)
    );

    fa fa_s4_c33_n15 (
        .a(stage4_col33[0]),
        .b(stage4_col33[1]),
        .c_in(stage4_col33[2]),
        .s(fa_s4_c33_n15_s),
        .c_out(fa_s4_c33_n15_c)
    );

    fa fa_s4_c34_n16 (
        .a(stage4_col34[0]),
        .b(stage4_col34[1]),
        .c_in(stage4_col34[2]),
        .s(fa_s4_c34_n16_s),
        .c_out(fa_s4_c34_n16_c)
    );

    fa fa_s4_c35_n17 (
        .a(stage4_col35[0]),
        .b(stage4_col35[1]),
        .c_in(stage4_col35[2]),
        .s(fa_s4_c35_n17_s),
        .c_out(fa_s4_c35_n17_c)
    );

    fa fa_s4_c36_n18 (
        .a(stage4_col36[0]),
        .b(stage4_col36[1]),
        .c_in(stage4_col36[2]),
        .s(fa_s4_c36_n18_s),
        .c_out(fa_s4_c36_n18_c)
    );

    fa fa_s4_c37_n19 (
        .a(stage4_col37[0]),
        .b(stage4_col37[1]),
        .c_in(stage4_col37[2]),
        .s(fa_s4_c37_n19_s),
        .c_out(fa_s4_c37_n19_c)
    );

    fa fa_s4_c38_n20 (
        .a(stage4_col38[0]),
        .b(stage4_col38[1]),
        .c_in(stage4_col38[2]),
        .s(fa_s4_c38_n20_s),
        .c_out(fa_s4_c38_n20_c)
    );

    fa fa_s4_c39_n21 (
        .a(stage4_col39[0]),
        .b(stage4_col39[1]),
        .c_in(stage4_col39[2]),
        .s(fa_s4_c39_n21_s),
        .c_out(fa_s4_c39_n21_c)
    );

    fa fa_s4_c40_n22 (
        .a(stage4_col40[0]),
        .b(stage4_col40[1]),
        .c_in(stage4_col40[2]),
        .s(fa_s4_c40_n22_s),
        .c_out(fa_s4_c40_n22_c)
    );

    fa fa_s4_c40_n23 (
        .a(stage4_col40[3]),
        .b(stage4_col40[4]),
        .c_in(stage4_col40[5]),
        .s(fa_s4_c40_n23_s),
        .c_out(fa_s4_c40_n23_c)
    );

    fa fa_s4_c41_n24 (
        .a(stage4_col41[0]),
        .b(stage4_col41[1]),
        .c_in(stage4_col41[2]),
        .s(fa_s4_c41_n24_s),
        .c_out(fa_s4_c41_n24_c)
    );

    fa fa_s4_c42_n25 (
        .a(stage4_col42[0]),
        .b(stage4_col42[1]),
        .c_in(stage4_col42[2]),
        .s(fa_s4_c42_n25_s),
        .c_out(fa_s4_c42_n25_c)
    );

    fa fa_s4_c43_n26 (
        .a(stage4_col43[0]),
        .b(stage4_col43[1]),
        .c_in(stage4_col43[2]),
        .s(fa_s4_c43_n26_s),
        .c_out(fa_s4_c43_n26_c)
    );

    fa fa_s4_c44_n27 (
        .a(stage4_col44[0]),
        .b(stage4_col44[1]),
        .c_in(stage4_col44[2]),
        .s(fa_s4_c44_n27_s),
        .c_out(fa_s4_c44_n27_c)
    );

    fa fa_s4_c45_n28 (
        .a(stage4_col45[0]),
        .b(stage4_col45[1]),
        .c_in(stage4_col45[2]),
        .s(fa_s4_c45_n28_s),
        .c_out(fa_s4_c45_n28_c)
    );

    fa fa_s4_c46_n29 (
        .a(stage4_col46[0]),
        .b(stage4_col46[1]),
        .c_in(stage4_col46[2]),
        .s(fa_s4_c46_n29_s),
        .c_out(fa_s4_c46_n29_c)
    );

    fa fa_s4_c47_n30 (
        .a(stage4_col47[0]),
        .b(stage4_col47[1]),
        .c_in(stage4_col47[2]),
        .s(fa_s4_c47_n30_s),
        .c_out(fa_s4_c47_n30_c)
    );

    fa fa_s4_c47_n31 (
        .a(stage4_col47[3]),
        .b(stage4_col47[4]),
        .c_in(stage4_col47[5]),
        .s(fa_s4_c47_n31_s),
        .c_out(fa_s4_c47_n31_c)
    );

    fa fa_s4_c48_n32 (
        .a(stage4_col48[0]),
        .b(stage4_col48[1]),
        .c_in(stage4_col48[2]),
        .s(fa_s4_c48_n32_s),
        .c_out(fa_s4_c48_n32_c)
    );

    fa fa_s4_c48_n33 (
        .a(stage4_col48[3]),
        .b(stage4_col48[4]),
        .c_in(stage4_col48[5]),
        .s(fa_s4_c48_n33_s),
        .c_out(fa_s4_c48_n33_c)
    );

    fa fa_s4_c49_n34 (
        .a(stage4_col49[0]),
        .b(stage4_col49[1]),
        .c_in(stage4_col49[2]),
        .s(fa_s4_c49_n34_s),
        .c_out(fa_s4_c49_n34_c)
    );

    fa fa_s4_c49_n35 (
        .a(stage4_col49[3]),
        .b(stage4_col49[4]),
        .c_in(stage4_col49[5]),
        .s(fa_s4_c49_n35_s),
        .c_out(fa_s4_c49_n35_c)
    );

    fa fa_s4_c50_n36 (
        .a(stage4_col50[0]),
        .b(stage4_col50[1]),
        .c_in(stage4_col50[2]),
        .s(fa_s4_c50_n36_s),
        .c_out(fa_s4_c50_n36_c)
    );

    fa fa_s4_c50_n37 (
        .a(stage4_col50[3]),
        .b(stage4_col50[4]),
        .c_in(stage4_col50[5]),
        .s(fa_s4_c50_n37_s),
        .c_out(fa_s4_c50_n37_c)
    );

    fa fa_s4_c51_n38 (
        .a(stage4_col51[0]),
        .b(stage4_col51[1]),
        .c_in(stage4_col51[2]),
        .s(fa_s4_c51_n38_s),
        .c_out(fa_s4_c51_n38_c)
    );

    fa fa_s4_c51_n39 (
        .a(stage4_col51[3]),
        .b(stage4_col51[4]),
        .c_in(stage4_col51[5]),
        .s(fa_s4_c51_n39_s),
        .c_out(fa_s4_c51_n39_c)
    );

    fa fa_s4_c52_n40 (
        .a(stage4_col52[0]),
        .b(stage4_col52[1]),
        .c_in(stage4_col52[2]),
        .s(fa_s4_c52_n40_s),
        .c_out(fa_s4_c52_n40_c)
    );

    fa fa_s4_c52_n41 (
        .a(stage4_col52[3]),
        .b(stage4_col52[4]),
        .c_in(stage4_col52[5]),
        .s(fa_s4_c52_n41_s),
        .c_out(fa_s4_c52_n41_c)
    );

    fa fa_s4_c53_n42 (
        .a(stage4_col53[0]),
        .b(stage4_col53[1]),
        .c_in(stage4_col53[2]),
        .s(fa_s4_c53_n42_s),
        .c_out(fa_s4_c53_n42_c)
    );

    fa fa_s4_c53_n43 (
        .a(stage4_col53[3]),
        .b(stage4_col53[4]),
        .c_in(stage4_col53[5]),
        .s(fa_s4_c53_n43_s),
        .c_out(fa_s4_c53_n43_c)
    );

    fa fa_s4_c54_n44 (
        .a(stage4_col54[0]),
        .b(stage4_col54[1]),
        .c_in(stage4_col54[2]),
        .s(fa_s4_c54_n44_s),
        .c_out(fa_s4_c54_n44_c)
    );

    fa fa_s4_c54_n45 (
        .a(stage4_col54[3]),
        .b(stage4_col54[4]),
        .c_in(stage4_col54[5]),
        .s(fa_s4_c54_n45_s),
        .c_out(fa_s4_c54_n45_c)
    );

    fa fa_s4_c55_n46 (
        .a(stage4_col55[0]),
        .b(stage4_col55[1]),
        .c_in(stage4_col55[2]),
        .s(fa_s4_c55_n46_s),
        .c_out(fa_s4_c55_n46_c)
    );

    fa fa_s4_c55_n47 (
        .a(stage4_col55[3]),
        .b(stage4_col55[4]),
        .c_in(stage4_col55[5]),
        .s(fa_s4_c55_n47_s),
        .c_out(fa_s4_c55_n47_c)
    );

    fa fa_s4_c56_n48 (
        .a(stage4_col56[0]),
        .b(stage4_col56[1]),
        .c_in(stage4_col56[2]),
        .s(fa_s4_c56_n48_s),
        .c_out(fa_s4_c56_n48_c)
    );

    fa fa_s4_c56_n49 (
        .a(stage4_col56[3]),
        .b(stage4_col56[4]),
        .c_in(stage4_col56[5]),
        .s(fa_s4_c56_n49_s),
        .c_out(fa_s4_c56_n49_c)
    );

    fa fa_s4_c57_n50 (
        .a(stage4_col57[0]),
        .b(stage4_col57[1]),
        .c_in(stage4_col57[2]),
        .s(fa_s4_c57_n50_s),
        .c_out(fa_s4_c57_n50_c)
    );

    fa fa_s4_c57_n51 (
        .a(stage4_col57[3]),
        .b(stage4_col57[4]),
        .c_in(stage4_col57[5]),
        .s(fa_s4_c57_n51_s),
        .c_out(fa_s4_c57_n51_c)
    );

    fa fa_s4_c58_n52 (
        .a(stage4_col58[0]),
        .b(stage4_col58[1]),
        .c_in(stage4_col58[2]),
        .s(fa_s4_c58_n52_s),
        .c_out(fa_s4_c58_n52_c)
    );

    fa fa_s4_c58_n53 (
        .a(stage4_col58[3]),
        .b(stage4_col58[4]),
        .c_in(stage4_col58[5]),
        .s(fa_s4_c58_n53_s),
        .c_out(fa_s4_c58_n53_c)
    );

    fa fa_s4_c59_n54 (
        .a(stage4_col59[0]),
        .b(stage4_col59[1]),
        .c_in(stage4_col59[2]),
        .s(fa_s4_c59_n54_s),
        .c_out(fa_s4_c59_n54_c)
    );

    fa fa_s4_c59_n55 (
        .a(stage4_col59[3]),
        .b(stage4_col59[4]),
        .c_in(stage4_col59[5]),
        .s(fa_s4_c59_n55_s),
        .c_out(fa_s4_c59_n55_c)
    );

    fa fa_s4_c60_n56 (
        .a(stage4_col60[0]),
        .b(stage4_col60[1]),
        .c_in(stage4_col60[2]),
        .s(fa_s4_c60_n56_s),
        .c_out(fa_s4_c60_n56_c)
    );

    fa fa_s4_c60_n57 (
        .a(stage4_col60[3]),
        .b(stage4_col60[4]),
        .c_in(stage4_col60[5]),
        .s(fa_s4_c60_n57_s),
        .c_out(fa_s4_c60_n57_c)
    );

    fa fa_s4_c61_n58 (
        .a(stage4_col61[0]),
        .b(stage4_col61[1]),
        .c_in(stage4_col61[2]),
        .s(fa_s4_c61_n58_s),
        .c_out(fa_s4_c61_n58_c)
    );

    fa fa_s4_c61_n59 (
        .a(stage4_col61[3]),
        .b(stage4_col61[4]),
        .c_in(stage4_col61[5]),
        .s(fa_s4_c61_n59_s),
        .c_out(fa_s4_c61_n59_c)
    );

    fa fa_s4_c62_n60 (
        .a(stage4_col62[0]),
        .b(stage4_col62[1]),
        .c_in(stage4_col62[2]),
        .s(fa_s4_c62_n60_s),
        .c_out(fa_s4_c62_n60_c)
    );

    fa fa_s4_c62_n61 (
        .a(stage4_col62[3]),
        .b(stage4_col62[4]),
        .c_in(stage4_col62[5]),
        .s(fa_s4_c62_n61_s),
        .c_out(fa_s4_c62_n61_c)
    );

    fa fa_s4_c63_n62 (
        .a(stage4_col63[0]),
        .b(stage4_col63[1]),
        .c_in(stage4_col63[2]),
        .s(fa_s4_c63_n62_s),
        .c_out(fa_s4_c63_n62_c)
    );

    fa fa_s4_c63_n63 (
        .a(stage4_col63[3]),
        .b(stage4_col63[4]),
        .c_in(stage4_col63[5]),
        .s(fa_s4_c63_n63_s),
        .c_out(fa_s4_c63_n63_c)
    );

    fa fa_s4_c64_n64 (
        .a(stage4_col64[0]),
        .b(stage4_col64[1]),
        .c_in(stage4_col64[2]),
        .s(fa_s4_c64_n64_s),
        .c_out(fa_s4_c64_n64_c)
    );

    fa fa_s4_c64_n65 (
        .a(stage4_col64[3]),
        .b(stage4_col64[4]),
        .c_in(stage4_col64[5]),
        .s(fa_s4_c64_n65_s),
        .c_out(fa_s4_c64_n65_c)
    );

    fa fa_s4_c65_n66 (
        .a(stage4_col65[0]),
        .b(stage4_col65[1]),
        .c_in(stage4_col65[2]),
        .s(fa_s4_c65_n66_s),
        .c_out(fa_s4_c65_n66_c)
    );

    fa fa_s4_c65_n67 (
        .a(stage4_col65[3]),
        .b(stage4_col65[4]),
        .c_in(stage4_col65[5]),
        .s(fa_s4_c65_n67_s),
        .c_out(fa_s4_c65_n67_c)
    );

    fa fa_s4_c66_n68 (
        .a(stage4_col66[0]),
        .b(stage4_col66[1]),
        .c_in(stage4_col66[2]),
        .s(fa_s4_c66_n68_s),
        .c_out(fa_s4_c66_n68_c)
    );

    fa fa_s4_c66_n69 (
        .a(stage4_col66[3]),
        .b(stage4_col66[4]),
        .c_in(stage4_col66[5]),
        .s(fa_s4_c66_n69_s),
        .c_out(fa_s4_c66_n69_c)
    );

    fa fa_s4_c67_n70 (
        .a(stage4_col67[0]),
        .b(stage4_col67[1]),
        .c_in(stage4_col67[2]),
        .s(fa_s4_c67_n70_s),
        .c_out(fa_s4_c67_n70_c)
    );

    fa fa_s4_c67_n71 (
        .a(stage4_col67[3]),
        .b(stage4_col67[4]),
        .c_in(stage4_col67[5]),
        .s(fa_s4_c67_n71_s),
        .c_out(fa_s4_c67_n71_c)
    );

    fa fa_s4_c68_n72 (
        .a(stage4_col68[0]),
        .b(stage4_col68[1]),
        .c_in(stage4_col68[2]),
        .s(fa_s4_c68_n72_s),
        .c_out(fa_s4_c68_n72_c)
    );

    fa fa_s4_c68_n73 (
        .a(stage4_col68[3]),
        .b(stage4_col68[4]),
        .c_in(stage4_col68[5]),
        .s(fa_s4_c68_n73_s),
        .c_out(fa_s4_c68_n73_c)
    );

    fa fa_s4_c69_n74 (
        .a(stage4_col69[0]),
        .b(stage4_col69[1]),
        .c_in(stage4_col69[2]),
        .s(fa_s4_c69_n74_s),
        .c_out(fa_s4_c69_n74_c)
    );

    fa fa_s4_c69_n75 (
        .a(stage4_col69[3]),
        .b(stage4_col69[4]),
        .c_in(stage4_col69[5]),
        .s(fa_s4_c69_n75_s),
        .c_out(fa_s4_c69_n75_c)
    );

    fa fa_s4_c70_n76 (
        .a(stage4_col70[0]),
        .b(stage4_col70[1]),
        .c_in(stage4_col70[2]),
        .s(fa_s4_c70_n76_s),
        .c_out(fa_s4_c70_n76_c)
    );

    fa fa_s4_c70_n77 (
        .a(stage4_col70[3]),
        .b(stage4_col70[4]),
        .c_in(stage4_col70[5]),
        .s(fa_s4_c70_n77_s),
        .c_out(fa_s4_c70_n77_c)
    );

    fa fa_s4_c71_n78 (
        .a(stage4_col71[0]),
        .b(stage4_col71[1]),
        .c_in(stage4_col71[2]),
        .s(fa_s4_c71_n78_s),
        .c_out(fa_s4_c71_n78_c)
    );

    fa fa_s4_c71_n79 (
        .a(stage4_col71[3]),
        .b(stage4_col71[4]),
        .c_in(stage4_col71[5]),
        .s(fa_s4_c71_n79_s),
        .c_out(fa_s4_c71_n79_c)
    );

    fa fa_s4_c72_n80 (
        .a(stage4_col72[0]),
        .b(stage4_col72[1]),
        .c_in(stage4_col72[2]),
        .s(fa_s4_c72_n80_s),
        .c_out(fa_s4_c72_n80_c)
    );

    fa fa_s4_c72_n81 (
        .a(stage4_col72[3]),
        .b(stage4_col72[4]),
        .c_in(stage4_col72[5]),
        .s(fa_s4_c72_n81_s),
        .c_out(fa_s4_c72_n81_c)
    );

    fa fa_s4_c73_n82 (
        .a(stage4_col73[0]),
        .b(stage4_col73[1]),
        .c_in(stage4_col73[2]),
        .s(fa_s4_c73_n82_s),
        .c_out(fa_s4_c73_n82_c)
    );

    fa fa_s4_c73_n83 (
        .a(stage4_col73[3]),
        .b(stage4_col73[4]),
        .c_in(stage4_col73[5]),
        .s(fa_s4_c73_n83_s),
        .c_out(fa_s4_c73_n83_c)
    );

    fa fa_s4_c74_n84 (
        .a(stage4_col74[0]),
        .b(stage4_col74[1]),
        .c_in(stage4_col74[2]),
        .s(fa_s4_c74_n84_s),
        .c_out(fa_s4_c74_n84_c)
    );

    fa fa_s4_c74_n85 (
        .a(stage4_col74[3]),
        .b(stage4_col74[4]),
        .c_in(stage4_col74[5]),
        .s(fa_s4_c74_n85_s),
        .c_out(fa_s4_c74_n85_c)
    );

    fa fa_s4_c75_n86 (
        .a(stage4_col75[0]),
        .b(stage4_col75[1]),
        .c_in(stage4_col75[2]),
        .s(fa_s4_c75_n86_s),
        .c_out(fa_s4_c75_n86_c)
    );

    fa fa_s4_c75_n87 (
        .a(stage4_col75[3]),
        .b(stage4_col75[4]),
        .c_in(stage4_col75[5]),
        .s(fa_s4_c75_n87_s),
        .c_out(fa_s4_c75_n87_c)
    );

    fa fa_s4_c76_n88 (
        .a(stage4_col76[0]),
        .b(stage4_col76[1]),
        .c_in(stage4_col76[2]),
        .s(fa_s4_c76_n88_s),
        .c_out(fa_s4_c76_n88_c)
    );

    fa fa_s4_c76_n89 (
        .a(stage4_col76[3]),
        .b(stage4_col76[4]),
        .c_in(stage4_col76[5]),
        .s(fa_s4_c76_n89_s),
        .c_out(fa_s4_c76_n89_c)
    );

    fa fa_s4_c77_n90 (
        .a(stage4_col77[0]),
        .b(stage4_col77[1]),
        .c_in(stage4_col77[2]),
        .s(fa_s4_c77_n90_s),
        .c_out(fa_s4_c77_n90_c)
    );

    fa fa_s4_c77_n91 (
        .a(stage4_col77[3]),
        .b(stage4_col77[4]),
        .c_in(stage4_col77[5]),
        .s(fa_s4_c77_n91_s),
        .c_out(fa_s4_c77_n91_c)
    );

    fa fa_s4_c78_n92 (
        .a(stage4_col78[0]),
        .b(stage4_col78[1]),
        .c_in(stage4_col78[2]),
        .s(fa_s4_c78_n92_s),
        .c_out(fa_s4_c78_n92_c)
    );

    fa fa_s4_c78_n93 (
        .a(stage4_col78[3]),
        .b(stage4_col78[4]),
        .c_in(stage4_col78[5]),
        .s(fa_s4_c78_n93_s),
        .c_out(fa_s4_c78_n93_c)
    );

    fa fa_s4_c79_n94 (
        .a(stage4_col79[0]),
        .b(stage4_col79[1]),
        .c_in(stage4_col79[2]),
        .s(fa_s4_c79_n94_s),
        .c_out(fa_s4_c79_n94_c)
    );

    fa fa_s4_c79_n95 (
        .a(stage4_col79[3]),
        .b(stage4_col79[4]),
        .c_in(stage4_col79[5]),
        .s(fa_s4_c79_n95_s),
        .c_out(fa_s4_c79_n95_c)
    );

    fa fa_s4_c80_n96 (
        .a(stage4_col80[0]),
        .b(stage4_col80[1]),
        .c_in(stage4_col80[2]),
        .s(fa_s4_c80_n96_s),
        .c_out(fa_s4_c80_n96_c)
    );

    fa fa_s4_c80_n97 (
        .a(stage4_col80[3]),
        .b(stage4_col80[4]),
        .c_in(stage4_col80[5]),
        .s(fa_s4_c80_n97_s),
        .c_out(fa_s4_c80_n97_c)
    );

    fa fa_s4_c81_n98 (
        .a(stage4_col81[0]),
        .b(stage4_col81[1]),
        .c_in(stage4_col81[2]),
        .s(fa_s4_c81_n98_s),
        .c_out(fa_s4_c81_n98_c)
    );

    fa fa_s4_c81_n99 (
        .a(stage4_col81[3]),
        .b(stage4_col81[4]),
        .c_in(stage4_col81[5]),
        .s(fa_s4_c81_n99_s),
        .c_out(fa_s4_c81_n99_c)
    );

    fa fa_s4_c82_n100 (
        .a(stage4_col82[0]),
        .b(stage4_col82[1]),
        .c_in(stage4_col82[2]),
        .s(fa_s4_c82_n100_s),
        .c_out(fa_s4_c82_n100_c)
    );

    fa fa_s4_c82_n101 (
        .a(stage4_col82[3]),
        .b(stage4_col82[4]),
        .c_in(stage4_col82[5]),
        .s(fa_s4_c82_n101_s),
        .c_out(fa_s4_c82_n101_c)
    );

    fa fa_s4_c83_n102 (
        .a(stage4_col83[0]),
        .b(stage4_col83[1]),
        .c_in(stage4_col83[2]),
        .s(fa_s4_c83_n102_s),
        .c_out(fa_s4_c83_n102_c)
    );

    fa fa_s4_c83_n103 (
        .a(stage4_col83[3]),
        .b(stage4_col83[4]),
        .c_in(stage4_col83[5]),
        .s(fa_s4_c83_n103_s),
        .c_out(fa_s4_c83_n103_c)
    );

    fa fa_s4_c84_n104 (
        .a(stage4_col84[0]),
        .b(stage4_col84[1]),
        .c_in(stage4_col84[2]),
        .s(fa_s4_c84_n104_s),
        .c_out(fa_s4_c84_n104_c)
    );

    fa fa_s4_c84_n105 (
        .a(stage4_col84[3]),
        .b(stage4_col84[4]),
        .c_in(stage4_col84[5]),
        .s(fa_s4_c84_n105_s),
        .c_out(fa_s4_c84_n105_c)
    );

    fa fa_s4_c85_n106 (
        .a(stage4_col85[0]),
        .b(stage4_col85[1]),
        .c_in(stage4_col85[2]),
        .s(fa_s4_c85_n106_s),
        .c_out(fa_s4_c85_n106_c)
    );

    fa fa_s4_c85_n107 (
        .a(stage4_col85[3]),
        .b(stage4_col85[4]),
        .c_in(stage4_col85[5]),
        .s(fa_s4_c85_n107_s),
        .c_out(fa_s4_c85_n107_c)
    );

    fa fa_s4_c86_n108 (
        .a(stage4_col86[0]),
        .b(stage4_col86[1]),
        .c_in(stage4_col86[2]),
        .s(fa_s4_c86_n108_s),
        .c_out(fa_s4_c86_n108_c)
    );

    fa fa_s4_c86_n109 (
        .a(stage4_col86[3]),
        .b(stage4_col86[4]),
        .c_in(stage4_col86[5]),
        .s(fa_s4_c86_n109_s),
        .c_out(fa_s4_c86_n109_c)
    );

    fa fa_s4_c87_n110 (
        .a(stage4_col87[0]),
        .b(stage4_col87[1]),
        .c_in(stage4_col87[2]),
        .s(fa_s4_c87_n110_s),
        .c_out(fa_s4_c87_n110_c)
    );

    fa fa_s4_c87_n111 (
        .a(stage4_col87[3]),
        .b(stage4_col87[4]),
        .c_in(stage4_col87[5]),
        .s(fa_s4_c87_n111_s),
        .c_out(fa_s4_c87_n111_c)
    );

    fa fa_s4_c88_n112 (
        .a(stage4_col88[0]),
        .b(stage4_col88[1]),
        .c_in(stage4_col88[2]),
        .s(fa_s4_c88_n112_s),
        .c_out(fa_s4_c88_n112_c)
    );

    fa fa_s4_c88_n113 (
        .a(stage4_col88[3]),
        .b(stage4_col88[4]),
        .c_in(stage4_col88[5]),
        .s(fa_s4_c88_n113_s),
        .c_out(fa_s4_c88_n113_c)
    );

    fa fa_s4_c89_n114 (
        .a(stage4_col89[0]),
        .b(stage4_col89[1]),
        .c_in(stage4_col89[2]),
        .s(fa_s4_c89_n114_s),
        .c_out(fa_s4_c89_n114_c)
    );

    fa fa_s4_c89_n115 (
        .a(stage4_col89[3]),
        .b(stage4_col89[4]),
        .c_in(stage4_col89[5]),
        .s(fa_s4_c89_n115_s),
        .c_out(fa_s4_c89_n115_c)
    );

    fa fa_s4_c90_n116 (
        .a(stage4_col90[0]),
        .b(stage4_col90[1]),
        .c_in(stage4_col90[2]),
        .s(fa_s4_c90_n116_s),
        .c_out(fa_s4_c90_n116_c)
    );

    fa fa_s4_c90_n117 (
        .a(stage4_col90[3]),
        .b(stage4_col90[4]),
        .c_in(stage4_col90[5]),
        .s(fa_s4_c90_n117_s),
        .c_out(fa_s4_c90_n117_c)
    );

    fa fa_s4_c91_n118 (
        .a(stage4_col91[0]),
        .b(stage4_col91[1]),
        .c_in(stage4_col91[2]),
        .s(fa_s4_c91_n118_s),
        .c_out(fa_s4_c91_n118_c)
    );

    fa fa_s4_c91_n119 (
        .a(stage4_col91[3]),
        .b(stage4_col91[4]),
        .c_in(stage4_col91[5]),
        .s(fa_s4_c91_n119_s),
        .c_out(fa_s4_c91_n119_c)
    );

    fa fa_s4_c92_n120 (
        .a(stage4_col92[0]),
        .b(stage4_col92[1]),
        .c_in(stage4_col92[2]),
        .s(fa_s4_c92_n120_s),
        .c_out(fa_s4_c92_n120_c)
    );

    fa fa_s4_c92_n121 (
        .a(stage4_col92[3]),
        .b(stage4_col92[4]),
        .c_in(stage4_col92[5]),
        .s(fa_s4_c92_n121_s),
        .c_out(fa_s4_c92_n121_c)
    );

    fa fa_s4_c93_n122 (
        .a(stage4_col93[0]),
        .b(stage4_col93[1]),
        .c_in(stage4_col93[2]),
        .s(fa_s4_c93_n122_s),
        .c_out(fa_s4_c93_n122_c)
    );

    fa fa_s4_c93_n123 (
        .a(stage4_col93[3]),
        .b(stage4_col93[4]),
        .c_in(stage4_col93[5]),
        .s(fa_s4_c93_n123_s),
        .c_out(fa_s4_c93_n123_c)
    );

    fa fa_s4_c94_n124 (
        .a(stage4_col94[0]),
        .b(stage4_col94[1]),
        .c_in(stage4_col94[2]),
        .s(fa_s4_c94_n124_s),
        .c_out(fa_s4_c94_n124_c)
    );

    fa fa_s4_c94_n125 (
        .a(stage4_col94[3]),
        .b(stage4_col94[4]),
        .c_in(stage4_col94[5]),
        .s(fa_s4_c94_n125_s),
        .c_out(fa_s4_c94_n125_c)
    );

    fa fa_s4_c95_n126 (
        .a(stage4_col95[0]),
        .b(stage4_col95[1]),
        .c_in(stage4_col95[2]),
        .s(fa_s4_c95_n126_s),
        .c_out(fa_s4_c95_n126_c)
    );

    fa fa_s4_c95_n127 (
        .a(stage4_col95[3]),
        .b(stage4_col95[4]),
        .c_in(stage4_col95[5]),
        .s(fa_s4_c95_n127_s),
        .c_out(fa_s4_c95_n127_c)
    );

    fa fa_s4_c96_n128 (
        .a(stage4_col96[0]),
        .b(stage4_col96[1]),
        .c_in(stage4_col96[2]),
        .s(fa_s4_c96_n128_s),
        .c_out(fa_s4_c96_n128_c)
    );

    fa fa_s4_c96_n129 (
        .a(stage4_col96[3]),
        .b(stage4_col96[4]),
        .c_in(stage4_col96[5]),
        .s(fa_s4_c96_n129_s),
        .c_out(fa_s4_c96_n129_c)
    );

    fa fa_s4_c97_n130 (
        .a(stage4_col97[0]),
        .b(stage4_col97[1]),
        .c_in(stage4_col97[2]),
        .s(fa_s4_c97_n130_s),
        .c_out(fa_s4_c97_n130_c)
    );

    fa fa_s4_c97_n131 (
        .a(stage4_col97[3]),
        .b(stage4_col97[4]),
        .c_in(stage4_col97[5]),
        .s(fa_s4_c97_n131_s),
        .c_out(fa_s4_c97_n131_c)
    );

    fa fa_s4_c98_n132 (
        .a(stage4_col98[0]),
        .b(stage4_col98[1]),
        .c_in(stage4_col98[2]),
        .s(fa_s4_c98_n132_s),
        .c_out(fa_s4_c98_n132_c)
    );

    fa fa_s4_c98_n133 (
        .a(stage4_col98[3]),
        .b(stage4_col98[4]),
        .c_in(stage4_col98[5]),
        .s(fa_s4_c98_n133_s),
        .c_out(fa_s4_c98_n133_c)
    );

    fa fa_s4_c99_n134 (
        .a(stage4_col99[0]),
        .b(stage4_col99[1]),
        .c_in(stage4_col99[2]),
        .s(fa_s4_c99_n134_s),
        .c_out(fa_s4_c99_n134_c)
    );

    fa fa_s4_c99_n135 (
        .a(stage4_col99[3]),
        .b(stage4_col99[4]),
        .c_in(stage4_col99[5]),
        .s(fa_s4_c99_n135_s),
        .c_out(fa_s4_c99_n135_c)
    );

    fa fa_s4_c100_n136 (
        .a(stage4_col100[0]),
        .b(stage4_col100[1]),
        .c_in(stage4_col100[2]),
        .s(fa_s4_c100_n136_s),
        .c_out(fa_s4_c100_n136_c)
    );

    fa fa_s4_c100_n137 (
        .a(stage4_col100[3]),
        .b(stage4_col100[4]),
        .c_in(stage4_col100[5]),
        .s(fa_s4_c100_n137_s),
        .c_out(fa_s4_c100_n137_c)
    );

    fa fa_s4_c101_n138 (
        .a(stage4_col101[0]),
        .b(stage4_col101[1]),
        .c_in(stage4_col101[2]),
        .s(fa_s4_c101_n138_s),
        .c_out(fa_s4_c101_n138_c)
    );

    fa fa_s4_c101_n139 (
        .a(stage4_col101[3]),
        .b(stage4_col101[4]),
        .c_in(stage4_col101[5]),
        .s(fa_s4_c101_n139_s),
        .c_out(fa_s4_c101_n139_c)
    );

    fa fa_s4_c102_n140 (
        .a(stage4_col102[0]),
        .b(stage4_col102[1]),
        .c_in(stage4_col102[2]),
        .s(fa_s4_c102_n140_s),
        .c_out(fa_s4_c102_n140_c)
    );

    fa fa_s4_c102_n141 (
        .a(stage4_col102[3]),
        .b(stage4_col102[4]),
        .c_in(stage4_col102[5]),
        .s(fa_s4_c102_n141_s),
        .c_out(fa_s4_c102_n141_c)
    );

    fa fa_s4_c103_n142 (
        .a(stage4_col103[0]),
        .b(stage4_col103[1]),
        .c_in(stage4_col103[2]),
        .s(fa_s4_c103_n142_s),
        .c_out(fa_s4_c103_n142_c)
    );

    fa fa_s4_c103_n143 (
        .a(stage4_col103[3]),
        .b(stage4_col103[4]),
        .c_in(stage4_col103[5]),
        .s(fa_s4_c103_n143_s),
        .c_out(fa_s4_c103_n143_c)
    );

    fa fa_s4_c104_n144 (
        .a(stage4_col104[0]),
        .b(stage4_col104[1]),
        .c_in(stage4_col104[2]),
        .s(fa_s4_c104_n144_s),
        .c_out(fa_s4_c104_n144_c)
    );

    fa fa_s4_c104_n145 (
        .a(stage4_col104[3]),
        .b(stage4_col104[4]),
        .c_in(stage4_col104[5]),
        .s(fa_s4_c104_n145_s),
        .c_out(fa_s4_c104_n145_c)
    );

    fa fa_s4_c105_n146 (
        .a(stage4_col105[0]),
        .b(stage4_col105[1]),
        .c_in(stage4_col105[2]),
        .s(fa_s4_c105_n146_s),
        .c_out(fa_s4_c105_n146_c)
    );

    fa fa_s4_c105_n147 (
        .a(stage4_col105[3]),
        .b(stage4_col105[4]),
        .c_in(stage4_col105[5]),
        .s(fa_s4_c105_n147_s),
        .c_out(fa_s4_c105_n147_c)
    );

    fa fa_s4_c106_n148 (
        .a(stage4_col106[0]),
        .b(stage4_col106[1]),
        .c_in(stage4_col106[2]),
        .s(fa_s4_c106_n148_s),
        .c_out(fa_s4_c106_n148_c)
    );

    fa fa_s4_c106_n149 (
        .a(stage4_col106[3]),
        .b(stage4_col106[4]),
        .c_in(stage4_col106[5]),
        .s(fa_s4_c106_n149_s),
        .c_out(fa_s4_c106_n149_c)
    );

    fa fa_s4_c107_n150 (
        .a(stage4_col107[0]),
        .b(stage4_col107[1]),
        .c_in(stage4_col107[2]),
        .s(fa_s4_c107_n150_s),
        .c_out(fa_s4_c107_n150_c)
    );

    fa fa_s4_c107_n151 (
        .a(stage4_col107[3]),
        .b(stage4_col107[4]),
        .c_in(stage4_col107[5]),
        .s(fa_s4_c107_n151_s),
        .c_out(fa_s4_c107_n151_c)
    );

    fa fa_s4_c108_n152 (
        .a(stage4_col108[0]),
        .b(stage4_col108[1]),
        .c_in(stage4_col108[2]),
        .s(fa_s4_c108_n152_s),
        .c_out(fa_s4_c108_n152_c)
    );

    fa fa_s4_c108_n153 (
        .a(stage4_col108[3]),
        .b(stage4_col108[4]),
        .c_in(stage4_col108[5]),
        .s(fa_s4_c108_n153_s),
        .c_out(fa_s4_c108_n153_c)
    );

    fa fa_s4_c109_n154 (
        .a(stage4_col109[0]),
        .b(stage4_col109[1]),
        .c_in(stage4_col109[2]),
        .s(fa_s4_c109_n154_s),
        .c_out(fa_s4_c109_n154_c)
    );

    fa fa_s4_c109_n155 (
        .a(stage4_col109[3]),
        .b(stage4_col109[4]),
        .c_in(stage4_col109[5]),
        .s(fa_s4_c109_n155_s),
        .c_out(fa_s4_c109_n155_c)
    );

    fa fa_s4_c110_n156 (
        .a(stage4_col110[0]),
        .b(stage4_col110[1]),
        .c_in(stage4_col110[2]),
        .s(fa_s4_c110_n156_s),
        .c_out(fa_s4_c110_n156_c)
    );

    fa fa_s4_c110_n157 (
        .a(stage4_col110[3]),
        .b(stage4_col110[4]),
        .c_in(stage4_col110[5]),
        .s(fa_s4_c110_n157_s),
        .c_out(fa_s4_c110_n157_c)
    );

    fa fa_s4_c111_n158 (
        .a(stage4_col111[0]),
        .b(stage4_col111[1]),
        .c_in(stage4_col111[2]),
        .s(fa_s4_c111_n158_s),
        .c_out(fa_s4_c111_n158_c)
    );

    fa fa_s4_c111_n159 (
        .a(stage4_col111[3]),
        .b(stage4_col111[4]),
        .c_in(stage4_col111[5]),
        .s(fa_s4_c111_n159_s),
        .c_out(fa_s4_c111_n159_c)
    );

    fa fa_s4_c112_n160 (
        .a(stage4_col112[0]),
        .b(stage4_col112[1]),
        .c_in(stage4_col112[2]),
        .s(fa_s4_c112_n160_s),
        .c_out(fa_s4_c112_n160_c)
    );

    fa fa_s4_c112_n161 (
        .a(stage4_col112[3]),
        .b(stage4_col112[4]),
        .c_in(stage4_col112[5]),
        .s(fa_s4_c112_n161_s),
        .c_out(fa_s4_c112_n161_c)
    );

    fa fa_s4_c113_n162 (
        .a(stage4_col113[0]),
        .b(stage4_col113[1]),
        .c_in(stage4_col113[2]),
        .s(fa_s4_c113_n162_s),
        .c_out(fa_s4_c113_n162_c)
    );

    fa fa_s4_c113_n163 (
        .a(stage4_col113[3]),
        .b(stage4_col113[4]),
        .c_in(stage4_col113[5]),
        .s(fa_s4_c113_n163_s),
        .c_out(fa_s4_c113_n163_c)
    );

    fa fa_s4_c114_n164 (
        .a(stage4_col114[0]),
        .b(stage4_col114[1]),
        .c_in(stage4_col114[2]),
        .s(fa_s4_c114_n164_s),
        .c_out(fa_s4_c114_n164_c)
    );

    fa fa_s4_c114_n165 (
        .a(stage4_col114[3]),
        .b(stage4_col114[4]),
        .c_in(stage4_col114[5]),
        .s(fa_s4_c114_n165_s),
        .c_out(fa_s4_c114_n165_c)
    );

    fa fa_s4_c115_n166 (
        .a(stage4_col115[0]),
        .b(stage4_col115[1]),
        .c_in(stage4_col115[2]),
        .s(fa_s4_c115_n166_s),
        .c_out(fa_s4_c115_n166_c)
    );

    fa fa_s4_c115_n167 (
        .a(stage4_col115[3]),
        .b(stage4_col115[4]),
        .c_in(stage4_col115[5]),
        .s(fa_s4_c115_n167_s),
        .c_out(fa_s4_c115_n167_c)
    );

    fa fa_s4_c116_n168 (
        .a(stage4_col116[0]),
        .b(stage4_col116[1]),
        .c_in(stage4_col116[2]),
        .s(fa_s4_c116_n168_s),
        .c_out(fa_s4_c116_n168_c)
    );

    fa fa_s4_c116_n169 (
        .a(stage4_col116[3]),
        .b(stage4_col116[4]),
        .c_in(stage4_col116[5]),
        .s(fa_s4_c116_n169_s),
        .c_out(fa_s4_c116_n169_c)
    );

    fa fa_s4_c117_n170 (
        .a(stage4_col117[0]),
        .b(stage4_col117[1]),
        .c_in(stage4_col117[2]),
        .s(fa_s4_c117_n170_s),
        .c_out(fa_s4_c117_n170_c)
    );

    fa fa_s4_c117_n171 (
        .a(stage4_col117[3]),
        .b(stage4_col117[4]),
        .c_in(stage4_col117[5]),
        .s(fa_s4_c117_n171_s),
        .c_out(fa_s4_c117_n171_c)
    );

    fa fa_s4_c118_n172 (
        .a(stage4_col118[0]),
        .b(stage4_col118[1]),
        .c_in(stage4_col118[2]),
        .s(fa_s4_c118_n172_s),
        .c_out(fa_s4_c118_n172_c)
    );

    fa fa_s4_c118_n173 (
        .a(stage4_col118[3]),
        .b(stage4_col118[4]),
        .c_in(stage4_col118[5]),
        .s(fa_s4_c118_n173_s),
        .c_out(fa_s4_c118_n173_c)
    );

    fa fa_s4_c119_n174 (
        .a(stage4_col119[0]),
        .b(stage4_col119[1]),
        .c_in(stage4_col119[2]),
        .s(fa_s4_c119_n174_s),
        .c_out(fa_s4_c119_n174_c)
    );

    fa fa_s4_c119_n175 (
        .a(stage4_col119[3]),
        .b(stage4_col119[4]),
        .c_in(stage4_col119[5]),
        .s(fa_s4_c119_n175_s),
        .c_out(fa_s4_c119_n175_c)
    );

    fa fa_s4_c120_n176 (
        .a(stage4_col120[0]),
        .b(stage4_col120[1]),
        .c_in(stage4_col120[2]),
        .s(fa_s4_c120_n176_s),
        .c_out(fa_s4_c120_n176_c)
    );

    fa fa_s4_c120_n177 (
        .a(stage4_col120[3]),
        .b(stage4_col120[4]),
        .c_in(stage4_col120[5]),
        .s(fa_s4_c120_n177_s),
        .c_out(fa_s4_c120_n177_c)
    );

    fa fa_s4_c121_n178 (
        .a(stage4_col121[0]),
        .b(stage4_col121[1]),
        .c_in(stage4_col121[2]),
        .s(fa_s4_c121_n178_s),
        .c_out(fa_s4_c121_n178_c)
    );

    fa fa_s4_c121_n179 (
        .a(stage4_col121[3]),
        .b(stage4_col121[4]),
        .c_in(stage4_col121[5]),
        .s(fa_s4_c121_n179_s),
        .c_out(fa_s4_c121_n179_c)
    );

    fa fa_s4_c122_n180 (
        .a(stage4_col122[0]),
        .b(stage4_col122[1]),
        .c_in(stage4_col122[2]),
        .s(fa_s4_c122_n180_s),
        .c_out(fa_s4_c122_n180_c)
    );

    fa fa_s4_c122_n181 (
        .a(stage4_col122[3]),
        .b(stage4_col122[4]),
        .c_in(stage4_col122[5]),
        .s(fa_s4_c122_n181_s),
        .c_out(fa_s4_c122_n181_c)
    );

    fa fa_s4_c123_n182 (
        .a(stage4_col123[0]),
        .b(stage4_col123[1]),
        .c_in(stage4_col123[2]),
        .s(fa_s4_c123_n182_s),
        .c_out(fa_s4_c123_n182_c)
    );

    fa fa_s4_c123_n183 (
        .a(stage4_col123[3]),
        .b(stage4_col123[4]),
        .c_in(stage4_col123[5]),
        .s(fa_s4_c123_n183_s),
        .c_out(fa_s4_c123_n183_c)
    );

    fa fa_s4_c124_n184 (
        .a(stage4_col124[0]),
        .b(stage4_col124[1]),
        .c_in(stage4_col124[2]),
        .s(fa_s4_c124_n184_s),
        .c_out(fa_s4_c124_n184_c)
    );

    fa fa_s4_c124_n185 (
        .a(stage4_col124[3]),
        .b(stage4_col124[4]),
        .c_in(stage4_col124[5]),
        .s(fa_s4_c124_n185_s),
        .c_out(fa_s4_c124_n185_c)
    );

    fa fa_s4_c125_n186 (
        .a(stage4_col125[0]),
        .b(stage4_col125[1]),
        .c_in(stage4_col125[2]),
        .s(fa_s4_c125_n186_s),
        .c_out(fa_s4_c125_n186_c)
    );

    fa fa_s4_c125_n187 (
        .a(stage4_col125[3]),
        .b(stage4_col125[4]),
        .c_in(stage4_col125[5]),
        .s(fa_s4_c125_n187_s),
        .c_out(fa_s4_c125_n187_c)
    );

    fa fa_s4_c126_n188 (
        .a(stage4_col126[0]),
        .b(stage4_col126[1]),
        .c_in(stage4_col126[2]),
        .s(fa_s4_c126_n188_s),
        .c_out(fa_s4_c126_n188_c)
    );

    fa fa_s4_c126_n189 (
        .a(stage4_col126[3]),
        .b(stage4_col126[4]),
        .c_in(stage4_col126[5]),
        .s(fa_s4_c126_n189_s),
        .c_out(fa_s4_c126_n189_c)
    );

    ha ha_s4_c4_n0 (
        .a(stage4_col4[0]),
        .b(stage4_col4[1]),
        .s(ha_s4_c4_n0_s),
        .c_out(ha_s4_c4_n0_c)
    );

    // Map to Stage 5 columns
    generate
        if (PIPE) begin : gen_stage5_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage5_col0[0] <= 1'b0;
                    stage5_col1[0] <= 1'b0;
                    stage5_col2[0] <= 1'b0;
                    stage5_col3[0] <= 1'b0;
                    stage5_col4[0] <= 1'b0;
                    stage5_col5[0] <= 1'b0;
                    stage5_col5[1] <= 1'b0;
                    stage5_col6[0] <= 1'b0;
                    stage5_col7[0] <= 1'b0;
                    stage5_col7[1] <= 1'b0;
                    stage5_col7[2] <= 1'b0;
                    stage5_col8[0] <= 1'b0;
                    stage5_col8[1] <= 1'b0;
                    stage5_col9[0] <= 1'b0;
                    stage5_col9[1] <= 1'b0;
                    stage5_col10[0] <= 1'b0;
                    stage5_col10[1] <= 1'b0;
                    stage5_col11[0] <= 1'b0;
                    stage5_col11[1] <= 1'b0;
                    stage5_col12[0] <= 1'b0;
                    stage5_col12[1] <= 1'b0;
                    stage5_col13[0] <= 1'b0;
                    stage5_col13[1] <= 1'b0;
                    stage5_col14[0] <= 1'b0;
                    stage5_col14[1] <= 1'b0;
                    stage5_col15[0] <= 1'b0;
                    stage5_col15[1] <= 1'b0;
                    stage5_col16[0] <= 1'b0;
                    stage5_col16[1] <= 1'b0;
                    stage5_col17[0] <= 1'b0;
                    stage5_col17[1] <= 1'b0;
                    stage5_col18[0] <= 1'b0;
                    stage5_col18[1] <= 1'b0;
                    stage5_col19[0] <= 1'b0;
                    stage5_col19[1] <= 1'b0;
                    stage5_col20[0] <= 1'b0;
                    stage5_col20[1] <= 1'b0;
                    stage5_col21[0] <= 1'b0;
                    stage5_col21[1] <= 1'b0;
                    stage5_col22[0] <= 1'b0;
                    stage5_col22[1] <= 1'b0;
                    stage5_col23[0] <= 1'b0;
                    stage5_col23[1] <= 1'b0;
                    stage5_col24[0] <= 1'b0;
                    stage5_col24[1] <= 1'b0;
                    stage5_col25[0] <= 1'b0;
                    stage5_col25[1] <= 1'b0;
                    stage5_col26[0] <= 1'b0;
                    stage5_col26[1] <= 1'b0;
                    stage5_col27[0] <= 1'b0;
                    stage5_col27[1] <= 1'b0;
                    stage5_col28[0] <= 1'b0;
                    stage5_col28[1] <= 1'b0;
                    stage5_col28[2] <= 1'b0;
                    stage5_col28[3] <= 1'b0;
                    stage5_col29[0] <= 1'b0;
                    stage5_col29[1] <= 1'b0;
                    stage5_col29[2] <= 1'b0;
                    stage5_col30[0] <= 1'b0;
                    stage5_col30[1] <= 1'b0;
                    stage5_col30[2] <= 1'b0;
                    stage5_col31[0] <= 1'b0;
                    stage5_col31[1] <= 1'b0;
                    stage5_col31[2] <= 1'b0;
                    stage5_col32[0] <= 1'b0;
                    stage5_col32[1] <= 1'b0;
                    stage5_col32[2] <= 1'b0;
                    stage5_col33[0] <= 1'b0;
                    stage5_col33[1] <= 1'b0;
                    stage5_col33[2] <= 1'b0;
                    stage5_col34[0] <= 1'b0;
                    stage5_col34[1] <= 1'b0;
                    stage5_col34[2] <= 1'b0;
                    stage5_col35[0] <= 1'b0;
                    stage5_col35[1] <= 1'b0;
                    stage5_col35[2] <= 1'b0;
                    stage5_col36[0] <= 1'b0;
                    stage5_col36[1] <= 1'b0;
                    stage5_col36[2] <= 1'b0;
                    stage5_col37[0] <= 1'b0;
                    stage5_col37[1] <= 1'b0;
                    stage5_col37[2] <= 1'b0;
                    stage5_col38[0] <= 1'b0;
                    stage5_col38[1] <= 1'b0;
                    stage5_col38[2] <= 1'b0;
                    stage5_col39[0] <= 1'b0;
                    stage5_col39[1] <= 1'b0;
                    stage5_col39[2] <= 1'b0;
                    stage5_col40[0] <= 1'b0;
                    stage5_col40[1] <= 1'b0;
                    stage5_col40[2] <= 1'b0;
                    stage5_col41[0] <= 1'b0;
                    stage5_col41[1] <= 1'b0;
                    stage5_col41[2] <= 1'b0;
                    stage5_col41[3] <= 1'b0;
                    stage5_col41[4] <= 1'b0;
                    stage5_col42[0] <= 1'b0;
                    stage5_col42[1] <= 1'b0;
                    stage5_col42[2] <= 1'b0;
                    stage5_col42[3] <= 1'b0;
                    stage5_col43[0] <= 1'b0;
                    stage5_col43[1] <= 1'b0;
                    stage5_col43[2] <= 1'b0;
                    stage5_col43[3] <= 1'b0;
                    stage5_col44[0] <= 1'b0;
                    stage5_col44[1] <= 1'b0;
                    stage5_col44[2] <= 1'b0;
                    stage5_col44[3] <= 1'b0;
                    stage5_col45[0] <= 1'b0;
                    stage5_col45[1] <= 1'b0;
                    stage5_col45[2] <= 1'b0;
                    stage5_col45[3] <= 1'b0;
                    stage5_col46[0] <= 1'b0;
                    stage5_col46[1] <= 1'b0;
                    stage5_col46[2] <= 1'b0;
                    stage5_col46[3] <= 1'b0;
                    stage5_col47[0] <= 1'b0;
                    stage5_col47[1] <= 1'b0;
                    stage5_col47[2] <= 1'b0;
                    stage5_col47[3] <= 1'b0;
                    stage5_col48[0] <= 1'b0;
                    stage5_col48[1] <= 1'b0;
                    stage5_col48[2] <= 1'b0;
                    stage5_col48[3] <= 1'b0;
                    stage5_col49[0] <= 1'b0;
                    stage5_col49[1] <= 1'b0;
                    stage5_col49[2] <= 1'b0;
                    stage5_col49[3] <= 1'b0;
                    stage5_col50[0] <= 1'b0;
                    stage5_col50[1] <= 1'b0;
                    stage5_col50[2] <= 1'b0;
                    stage5_col50[3] <= 1'b0;
                    stage5_col51[0] <= 1'b0;
                    stage5_col51[1] <= 1'b0;
                    stage5_col51[2] <= 1'b0;
                    stage5_col51[3] <= 1'b0;
                    stage5_col52[0] <= 1'b0;
                    stage5_col52[1] <= 1'b0;
                    stage5_col52[2] <= 1'b0;
                    stage5_col52[3] <= 1'b0;
                    stage5_col53[0] <= 1'b0;
                    stage5_col53[1] <= 1'b0;
                    stage5_col53[2] <= 1'b0;
                    stage5_col53[3] <= 1'b0;
                    stage5_col54[0] <= 1'b0;
                    stage5_col54[1] <= 1'b0;
                    stage5_col54[2] <= 1'b0;
                    stage5_col54[3] <= 1'b0;
                    stage5_col55[0] <= 1'b0;
                    stage5_col55[1] <= 1'b0;
                    stage5_col55[2] <= 1'b0;
                    stage5_col55[3] <= 1'b0;
                    stage5_col56[0] <= 1'b0;
                    stage5_col56[1] <= 1'b0;
                    stage5_col56[2] <= 1'b0;
                    stage5_col56[3] <= 1'b0;
                    stage5_col57[0] <= 1'b0;
                    stage5_col57[1] <= 1'b0;
                    stage5_col57[2] <= 1'b0;
                    stage5_col57[3] <= 1'b0;
                    stage5_col58[0] <= 1'b0;
                    stage5_col58[1] <= 1'b0;
                    stage5_col58[2] <= 1'b0;
                    stage5_col58[3] <= 1'b0;
                    stage5_col59[0] <= 1'b0;
                    stage5_col59[1] <= 1'b0;
                    stage5_col59[2] <= 1'b0;
                    stage5_col59[3] <= 1'b0;
                    stage5_col59[4] <= 1'b0;
                    stage5_col59[5] <= 1'b0;
                    stage5_col60[0] <= 1'b0;
                    stage5_col60[1] <= 1'b0;
                    stage5_col60[2] <= 1'b0;
                    stage5_col60[3] <= 1'b0;
                    stage5_col60[4] <= 1'b0;
                    stage5_col61[0] <= 1'b0;
                    stage5_col61[1] <= 1'b0;
                    stage5_col61[2] <= 1'b0;
                    stage5_col61[3] <= 1'b0;
                    stage5_col61[4] <= 1'b0;
                    stage5_col62[0] <= 1'b0;
                    stage5_col62[1] <= 1'b0;
                    stage5_col62[2] <= 1'b0;
                    stage5_col62[3] <= 1'b0;
                    stage5_col62[4] <= 1'b0;
                    stage5_col63[0] <= 1'b0;
                    stage5_col63[1] <= 1'b0;
                    stage5_col63[2] <= 1'b0;
                    stage5_col63[3] <= 1'b0;
                    stage5_col63[4] <= 1'b0;
                    stage5_col64[0] <= 1'b0;
                    stage5_col64[1] <= 1'b0;
                    stage5_col64[2] <= 1'b0;
                    stage5_col64[3] <= 1'b0;
                    stage5_col64[4] <= 1'b0;
                    stage5_col64[5] <= 1'b0;
                    stage5_col65[0] <= 1'b0;
                    stage5_col65[1] <= 1'b0;
                    stage5_col65[2] <= 1'b0;
                    stage5_col65[3] <= 1'b0;
                    stage5_col65[4] <= 1'b0;
                    stage5_col66[0] <= 1'b0;
                    stage5_col66[1] <= 1'b0;
                    stage5_col66[2] <= 1'b0;
                    stage5_col66[3] <= 1'b0;
                    stage5_col66[4] <= 1'b0;
                    stage5_col66[5] <= 1'b0;
                    stage5_col67[0] <= 1'b0;
                    stage5_col67[1] <= 1'b0;
                    stage5_col67[2] <= 1'b0;
                    stage5_col67[3] <= 1'b0;
                    stage5_col67[4] <= 1'b0;
                    stage5_col68[0] <= 1'b0;
                    stage5_col68[1] <= 1'b0;
                    stage5_col68[2] <= 1'b0;
                    stage5_col68[3] <= 1'b0;
                    stage5_col68[4] <= 1'b0;
                    stage5_col68[5] <= 1'b0;
                    stage5_col69[0] <= 1'b0;
                    stage5_col69[1] <= 1'b0;
                    stage5_col69[2] <= 1'b0;
                    stage5_col69[3] <= 1'b0;
                    stage5_col69[4] <= 1'b0;
                    stage5_col70[0] <= 1'b0;
                    stage5_col70[1] <= 1'b0;
                    stage5_col70[2] <= 1'b0;
                    stage5_col70[3] <= 1'b0;
                    stage5_col70[4] <= 1'b0;
                    stage5_col70[5] <= 1'b0;
                    stage5_col71[0] <= 1'b0;
                    stage5_col71[1] <= 1'b0;
                    stage5_col71[2] <= 1'b0;
                    stage5_col71[3] <= 1'b0;
                    stage5_col71[4] <= 1'b0;
                    stage5_col72[0] <= 1'b0;
                    stage5_col72[1] <= 1'b0;
                    stage5_col72[2] <= 1'b0;
                    stage5_col72[3] <= 1'b0;
                    stage5_col72[4] <= 1'b0;
                    stage5_col72[5] <= 1'b0;
                    stage5_col73[0] <= 1'b0;
                    stage5_col73[1] <= 1'b0;
                    stage5_col73[2] <= 1'b0;
                    stage5_col73[3] <= 1'b0;
                    stage5_col73[4] <= 1'b0;
                    stage5_col74[0] <= 1'b0;
                    stage5_col74[1] <= 1'b0;
                    stage5_col74[2] <= 1'b0;
                    stage5_col74[3] <= 1'b0;
                    stage5_col74[4] <= 1'b0;
                    stage5_col74[5] <= 1'b0;
                    stage5_col75[0] <= 1'b0;
                    stage5_col75[1] <= 1'b0;
                    stage5_col75[2] <= 1'b0;
                    stage5_col75[3] <= 1'b0;
                    stage5_col75[4] <= 1'b0;
                    stage5_col76[0] <= 1'b0;
                    stage5_col76[1] <= 1'b0;
                    stage5_col76[2] <= 1'b0;
                    stage5_col76[3] <= 1'b0;
                    stage5_col76[4] <= 1'b0;
                    stage5_col76[5] <= 1'b0;
                    stage5_col77[0] <= 1'b0;
                    stage5_col77[1] <= 1'b0;
                    stage5_col77[2] <= 1'b0;
                    stage5_col77[3] <= 1'b0;
                    stage5_col77[4] <= 1'b0;
                    stage5_col78[0] <= 1'b0;
                    stage5_col78[1] <= 1'b0;
                    stage5_col78[2] <= 1'b0;
                    stage5_col78[3] <= 1'b0;
                    stage5_col78[4] <= 1'b0;
                    stage5_col78[5] <= 1'b0;
                    stage5_col79[0] <= 1'b0;
                    stage5_col79[1] <= 1'b0;
                    stage5_col79[2] <= 1'b0;
                    stage5_col79[3] <= 1'b0;
                    stage5_col79[4] <= 1'b0;
                    stage5_col80[0] <= 1'b0;
                    stage5_col80[1] <= 1'b0;
                    stage5_col80[2] <= 1'b0;
                    stage5_col80[3] <= 1'b0;
                    stage5_col80[4] <= 1'b0;
                    stage5_col80[5] <= 1'b0;
                    stage5_col81[0] <= 1'b0;
                    stage5_col81[1] <= 1'b0;
                    stage5_col81[2] <= 1'b0;
                    stage5_col81[3] <= 1'b0;
                    stage5_col81[4] <= 1'b0;
                    stage5_col82[0] <= 1'b0;
                    stage5_col82[1] <= 1'b0;
                    stage5_col82[2] <= 1'b0;
                    stage5_col82[3] <= 1'b0;
                    stage5_col82[4] <= 1'b0;
                    stage5_col82[5] <= 1'b0;
                    stage5_col83[0] <= 1'b0;
                    stage5_col83[1] <= 1'b0;
                    stage5_col83[2] <= 1'b0;
                    stage5_col83[3] <= 1'b0;
                    stage5_col83[4] <= 1'b0;
                    stage5_col84[0] <= 1'b0;
                    stage5_col84[1] <= 1'b0;
                    stage5_col84[2] <= 1'b0;
                    stage5_col84[3] <= 1'b0;
                    stage5_col84[4] <= 1'b0;
                    stage5_col84[5] <= 1'b0;
                    stage5_col85[0] <= 1'b0;
                    stage5_col85[1] <= 1'b0;
                    stage5_col85[2] <= 1'b0;
                    stage5_col85[3] <= 1'b0;
                    stage5_col85[4] <= 1'b0;
                    stage5_col86[0] <= 1'b0;
                    stage5_col86[1] <= 1'b0;
                    stage5_col86[2] <= 1'b0;
                    stage5_col86[3] <= 1'b0;
                    stage5_col86[4] <= 1'b0;
                    stage5_col86[5] <= 1'b0;
                    stage5_col87[0] <= 1'b0;
                    stage5_col87[1] <= 1'b0;
                    stage5_col87[2] <= 1'b0;
                    stage5_col87[3] <= 1'b0;
                    stage5_col87[4] <= 1'b0;
                    stage5_col88[0] <= 1'b0;
                    stage5_col88[1] <= 1'b0;
                    stage5_col88[2] <= 1'b0;
                    stage5_col88[3] <= 1'b0;
                    stage5_col88[4] <= 1'b0;
                    stage5_col88[5] <= 1'b0;
                    stage5_col89[0] <= 1'b0;
                    stage5_col89[1] <= 1'b0;
                    stage5_col89[2] <= 1'b0;
                    stage5_col89[3] <= 1'b0;
                    stage5_col89[4] <= 1'b0;
                    stage5_col90[0] <= 1'b0;
                    stage5_col90[1] <= 1'b0;
                    stage5_col90[2] <= 1'b0;
                    stage5_col90[3] <= 1'b0;
                    stage5_col90[4] <= 1'b0;
                    stage5_col90[5] <= 1'b0;
                    stage5_col91[0] <= 1'b0;
                    stage5_col91[1] <= 1'b0;
                    stage5_col91[2] <= 1'b0;
                    stage5_col91[3] <= 1'b0;
                    stage5_col91[4] <= 1'b0;
                    stage5_col92[0] <= 1'b0;
                    stage5_col92[1] <= 1'b0;
                    stage5_col92[2] <= 1'b0;
                    stage5_col92[3] <= 1'b0;
                    stage5_col92[4] <= 1'b0;
                    stage5_col92[5] <= 1'b0;
                    stage5_col93[0] <= 1'b0;
                    stage5_col93[1] <= 1'b0;
                    stage5_col93[2] <= 1'b0;
                    stage5_col93[3] <= 1'b0;
                    stage5_col93[4] <= 1'b0;
                    stage5_col94[0] <= 1'b0;
                    stage5_col94[1] <= 1'b0;
                    stage5_col94[2] <= 1'b0;
                    stage5_col94[3] <= 1'b0;
                    stage5_col94[4] <= 1'b0;
                    stage5_col94[5] <= 1'b0;
                    stage5_col95[0] <= 1'b0;
                    stage5_col95[1] <= 1'b0;
                    stage5_col95[2] <= 1'b0;
                    stage5_col95[3] <= 1'b0;
                    stage5_col95[4] <= 1'b0;
                    stage5_col96[0] <= 1'b0;
                    stage5_col96[1] <= 1'b0;
                    stage5_col96[2] <= 1'b0;
                    stage5_col96[3] <= 1'b0;
                    stage5_col96[4] <= 1'b0;
                    stage5_col96[5] <= 1'b0;
                    stage5_col97[0] <= 1'b0;
                    stage5_col97[1] <= 1'b0;
                    stage5_col97[2] <= 1'b0;
                    stage5_col97[3] <= 1'b0;
                    stage5_col97[4] <= 1'b0;
                    stage5_col98[0] <= 1'b0;
                    stage5_col98[1] <= 1'b0;
                    stage5_col98[2] <= 1'b0;
                    stage5_col98[3] <= 1'b0;
                    stage5_col98[4] <= 1'b0;
                    stage5_col98[5] <= 1'b0;
                    stage5_col99[0] <= 1'b0;
                    stage5_col99[1] <= 1'b0;
                    stage5_col99[2] <= 1'b0;
                    stage5_col99[3] <= 1'b0;
                    stage5_col99[4] <= 1'b0;
                    stage5_col100[0] <= 1'b0;
                    stage5_col100[1] <= 1'b0;
                    stage5_col100[2] <= 1'b0;
                    stage5_col100[3] <= 1'b0;
                    stage5_col100[4] <= 1'b0;
                    stage5_col100[5] <= 1'b0;
                    stage5_col101[0] <= 1'b0;
                    stage5_col101[1] <= 1'b0;
                    stage5_col101[2] <= 1'b0;
                    stage5_col101[3] <= 1'b0;
                    stage5_col101[4] <= 1'b0;
                    stage5_col102[0] <= 1'b0;
                    stage5_col102[1] <= 1'b0;
                    stage5_col102[2] <= 1'b0;
                    stage5_col102[3] <= 1'b0;
                    stage5_col102[4] <= 1'b0;
                    stage5_col102[5] <= 1'b0;
                    stage5_col103[0] <= 1'b0;
                    stage5_col103[1] <= 1'b0;
                    stage5_col103[2] <= 1'b0;
                    stage5_col103[3] <= 1'b0;
                    stage5_col103[4] <= 1'b0;
                    stage5_col104[0] <= 1'b0;
                    stage5_col104[1] <= 1'b0;
                    stage5_col104[2] <= 1'b0;
                    stage5_col104[3] <= 1'b0;
                    stage5_col104[4] <= 1'b0;
                    stage5_col104[5] <= 1'b0;
                    stage5_col105[0] <= 1'b0;
                    stage5_col105[1] <= 1'b0;
                    stage5_col105[2] <= 1'b0;
                    stage5_col105[3] <= 1'b0;
                    stage5_col105[4] <= 1'b0;
                    stage5_col106[0] <= 1'b0;
                    stage5_col106[1] <= 1'b0;
                    stage5_col106[2] <= 1'b0;
                    stage5_col106[3] <= 1'b0;
                    stage5_col106[4] <= 1'b0;
                    stage5_col106[5] <= 1'b0;
                    stage5_col107[0] <= 1'b0;
                    stage5_col107[1] <= 1'b0;
                    stage5_col107[2] <= 1'b0;
                    stage5_col107[3] <= 1'b0;
                    stage5_col107[4] <= 1'b0;
                    stage5_col108[0] <= 1'b0;
                    stage5_col108[1] <= 1'b0;
                    stage5_col108[2] <= 1'b0;
                    stage5_col108[3] <= 1'b0;
                    stage5_col108[4] <= 1'b0;
                    stage5_col108[5] <= 1'b0;
                    stage5_col109[0] <= 1'b0;
                    stage5_col109[1] <= 1'b0;
                    stage5_col109[2] <= 1'b0;
                    stage5_col109[3] <= 1'b0;
                    stage5_col109[4] <= 1'b0;
                    stage5_col110[0] <= 1'b0;
                    stage5_col110[1] <= 1'b0;
                    stage5_col110[2] <= 1'b0;
                    stage5_col110[3] <= 1'b0;
                    stage5_col110[4] <= 1'b0;
                    stage5_col110[5] <= 1'b0;
                    stage5_col111[0] <= 1'b0;
                    stage5_col111[1] <= 1'b0;
                    stage5_col111[2] <= 1'b0;
                    stage5_col111[3] <= 1'b0;
                    stage5_col111[4] <= 1'b0;
                    stage5_col112[0] <= 1'b0;
                    stage5_col112[1] <= 1'b0;
                    stage5_col112[2] <= 1'b0;
                    stage5_col112[3] <= 1'b0;
                    stage5_col112[4] <= 1'b0;
                    stage5_col112[5] <= 1'b0;
                    stage5_col113[0] <= 1'b0;
                    stage5_col113[1] <= 1'b0;
                    stage5_col113[2] <= 1'b0;
                    stage5_col113[3] <= 1'b0;
                    stage5_col113[4] <= 1'b0;
                    stage5_col114[0] <= 1'b0;
                    stage5_col114[1] <= 1'b0;
                    stage5_col114[2] <= 1'b0;
                    stage5_col114[3] <= 1'b0;
                    stage5_col114[4] <= 1'b0;
                    stage5_col114[5] <= 1'b0;
                    stage5_col115[0] <= 1'b0;
                    stage5_col115[1] <= 1'b0;
                    stage5_col115[2] <= 1'b0;
                    stage5_col115[3] <= 1'b0;
                    stage5_col115[4] <= 1'b0;
                    stage5_col116[0] <= 1'b0;
                    stage5_col116[1] <= 1'b0;
                    stage5_col116[2] <= 1'b0;
                    stage5_col116[3] <= 1'b0;
                    stage5_col116[4] <= 1'b0;
                    stage5_col116[5] <= 1'b0;
                    stage5_col117[0] <= 1'b0;
                    stage5_col117[1] <= 1'b0;
                    stage5_col117[2] <= 1'b0;
                    stage5_col117[3] <= 1'b0;
                    stage5_col117[4] <= 1'b0;
                    stage5_col118[0] <= 1'b0;
                    stage5_col118[1] <= 1'b0;
                    stage5_col118[2] <= 1'b0;
                    stage5_col118[3] <= 1'b0;
                    stage5_col118[4] <= 1'b0;
                    stage5_col118[5] <= 1'b0;
                    stage5_col119[0] <= 1'b0;
                    stage5_col119[1] <= 1'b0;
                    stage5_col119[2] <= 1'b0;
                    stage5_col119[3] <= 1'b0;
                    stage5_col119[4] <= 1'b0;
                    stage5_col120[0] <= 1'b0;
                    stage5_col120[1] <= 1'b0;
                    stage5_col120[2] <= 1'b0;
                    stage5_col120[3] <= 1'b0;
                    stage5_col120[4] <= 1'b0;
                    stage5_col120[5] <= 1'b0;
                    stage5_col121[0] <= 1'b0;
                    stage5_col121[1] <= 1'b0;
                    stage5_col121[2] <= 1'b0;
                    stage5_col121[3] <= 1'b0;
                    stage5_col121[4] <= 1'b0;
                    stage5_col122[0] <= 1'b0;
                    stage5_col122[1] <= 1'b0;
                    stage5_col122[2] <= 1'b0;
                    stage5_col122[3] <= 1'b0;
                    stage5_col122[4] <= 1'b0;
                    stage5_col122[5] <= 1'b0;
                    stage5_col123[0] <= 1'b0;
                    stage5_col123[1] <= 1'b0;
                    stage5_col123[2] <= 1'b0;
                    stage5_col123[3] <= 1'b0;
                    stage5_col123[4] <= 1'b0;
                    stage5_col124[0] <= 1'b0;
                    stage5_col124[1] <= 1'b0;
                    stage5_col124[2] <= 1'b0;
                    stage5_col124[3] <= 1'b0;
                    stage5_col124[4] <= 1'b0;
                    stage5_col124[5] <= 1'b0;
                    stage5_col125[0] <= 1'b0;
                    stage5_col125[1] <= 1'b0;
                    stage5_col125[2] <= 1'b0;
                    stage5_col125[3] <= 1'b0;
                    stage5_col125[4] <= 1'b0;
                    stage5_col126[0] <= 1'b0;
                    stage5_col126[1] <= 1'b0;
                    stage5_col126[2] <= 1'b0;
                    stage5_col126[3] <= 1'b0;
                    stage5_col126[4] <= 1'b0;
                    stage5_col126[5] <= 1'b0;
                    stage5_col127[0] <= 1'b0;
                    stage5_col127[1] <= 1'b0;
                    stage5_col127[2] <= 1'b0;
                    stage5_col127[3] <= 1'b0;
                    stage5_col127[4] <= 1'b0;
                    stage5_col127[5] <= 1'b0;
                    stage5_col127[6] <= 1'b0;
                    stage5_col127[7] <= 1'b0;
                    stage5_col127[8] <= 1'b0;
                    stage5_col127[9] <= 1'b0;
                    stage5_col127[10] <= 1'b0;
                    stage5_col127[11] <= 1'b0;
                    stage5_col127[12] <= 1'b0;
                    stage5_col127[13] <= 1'b0;
                    stage5_col127[14] <= 1'b0;
                    stage5_col127[15] <= 1'b0;
                    stage5_col127[16] <= 1'b0;
                    stage5_col127[17] <= 1'b0;
                    stage5_col127[18] <= 1'b0;
                    stage5_col127[19] <= 1'b0;
                    stage5_col127[20] <= 1'b0;
                    stage5_col127[21] <= 1'b0;
                    stage5_col127[22] <= 1'b0;
                    stage5_col127[23] <= 1'b0;
                    stage5_col127[24] <= 1'b0;
                    stage5_col127[25] <= 1'b0;
                    stage5_col127[26] <= 1'b0;
                    stage5_col127[27] <= 1'b0;
                    stage5_col127[28] <= 1'b0;
                    stage5_col127[29] <= 1'b0;
                    stage5_col127[30] <= 1'b0;
                    stage5_col127[31] <= 1'b0;
                    stage5_col127[32] <= 1'b0;
                    stage5_col127[33] <= 1'b0;
                    stage5_col127[34] <= 1'b0;
                    stage5_col127[35] <= 1'b0;
                    stage5_col127[36] <= 1'b0;
                    stage5_col127[37] <= 1'b0;
                    stage5_col127[38] <= 1'b0;
                    stage5_col127[39] <= 1'b0;
                    stage5_col127[40] <= 1'b0;
                    stage5_col127[41] <= 1'b0;
                    stage5_col127[42] <= 1'b0;
                    stage5_col127[43] <= 1'b0;
                    stage5_col127[44] <= 1'b0;
                    stage5_col127[45] <= 1'b0;
                    stage5_col127[46] <= 1'b0;
                    stage5_col127[47] <= 1'b0;
                    stage5_col127[48] <= 1'b0;
                    stage5_col127[49] <= 1'b0;
                    stage5_col127[50] <= 1'b0;
                    stage5_col127[51] <= 1'b0;
                    stage5_col127[52] <= 1'b0;
                    stage5_col127[53] <= 1'b0;
                    stage5_col127[54] <= 1'b0;
                    stage5_col127[55] <= 1'b0;
                    stage5_col127[56] <= 1'b0;
                    stage5_col127[57] <= 1'b0;
                    stage5_col127[58] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage5_col0[0] <= stage4_col0[0];
                    stage5_col1[0] <= stage4_col1[0];
                    stage5_col2[0] <= stage4_col2[0];
                    stage5_col3[0] <= stage4_col3[0];
                    stage5_col4[0] <= ha_s4_c4_n0_s;
                    stage5_col5[0] <= ha_s4_c4_n0_c;
                    stage5_col5[1] <= stage4_col5[0];
                    stage5_col6[0] <= fa_s4_c6_n0_s;
                    stage5_col7[0] <= fa_s4_c6_n0_c;
                    stage5_col7[1] <= stage4_col7[0];
                    stage5_col7[2] <= stage4_col7[1];
                    stage5_col8[0] <= stage4_col8[0];
                    stage5_col8[1] <= stage4_col8[1];
                    stage5_col9[0] <= stage4_col9[0];
                    stage5_col9[1] <= stage4_col9[1];
                    stage5_col10[0] <= stage4_col10[0];
                    stage5_col10[1] <= stage4_col10[1];
                    stage5_col11[0] <= stage4_col11[0];
                    stage5_col11[1] <= stage4_col11[1];
                    stage5_col12[0] <= stage4_col12[0];
                    stage5_col12[1] <= stage4_col12[1];
                    stage5_col13[0] <= stage4_col13[0];
                    stage5_col13[1] <= stage4_col13[1];
                    stage5_col14[0] <= stage4_col14[0];
                    stage5_col14[1] <= stage4_col14[1];
                    stage5_col15[0] <= stage4_col15[0];
                    stage5_col15[1] <= stage4_col15[1];
                    stage5_col16[0] <= stage4_col16[0];
                    stage5_col16[1] <= stage4_col16[1];
                    stage5_col17[0] <= stage4_col17[0];
                    stage5_col17[1] <= stage4_col17[1];
                    stage5_col18[0] <= stage4_col18[0];
                    stage5_col18[1] <= stage4_col18[1];
                    stage5_col19[0] <= fa_s4_c19_n1_s;
                    stage5_col19[1] <= stage4_col19[3];
                    stage5_col20[0] <= fa_s4_c19_n1_c;
                    stage5_col20[1] <= fa_s4_c20_n2_s;
                    stage5_col21[0] <= fa_s4_c20_n2_c;
                    stage5_col21[1] <= fa_s4_c21_n3_s;
                    stage5_col22[0] <= fa_s4_c21_n3_c;
                    stage5_col22[1] <= fa_s4_c22_n4_s;
                    stage5_col23[0] <= fa_s4_c22_n4_c;
                    stage5_col23[1] <= fa_s4_c23_n5_s;
                    stage5_col24[0] <= fa_s4_c23_n5_c;
                    stage5_col24[1] <= fa_s4_c24_n6_s;
                    stage5_col25[0] <= fa_s4_c24_n6_c;
                    stage5_col25[1] <= fa_s4_c25_n7_s;
                    stage5_col26[0] <= fa_s4_c25_n7_c;
                    stage5_col26[1] <= fa_s4_c26_n8_s;
                    stage5_col27[0] <= fa_s4_c26_n8_c;
                    stage5_col27[1] <= fa_s4_c27_n9_s;
                    stage5_col28[0] <= fa_s4_c27_n9_c;
                    stage5_col28[1] <= fa_s4_c28_n10_s;
                    stage5_col28[2] <= stage4_col28[3];
                    stage5_col28[3] <= stage4_col28[4];
                    stage5_col29[0] <= fa_s4_c28_n10_c;
                    stage5_col29[1] <= fa_s4_c29_n11_s;
                    stage5_col29[2] <= stage4_col29[3];
                    stage5_col30[0] <= fa_s4_c29_n11_c;
                    stage5_col30[1] <= fa_s4_c30_n12_s;
                    stage5_col30[2] <= stage4_col30[3];
                    stage5_col31[0] <= fa_s4_c30_n12_c;
                    stage5_col31[1] <= fa_s4_c31_n13_s;
                    stage5_col31[2] <= stage4_col31[3];
                    stage5_col32[0] <= fa_s4_c31_n13_c;
                    stage5_col32[1] <= fa_s4_c32_n14_s;
                    stage5_col32[2] <= stage4_col32[3];
                    stage5_col33[0] <= fa_s4_c32_n14_c;
                    stage5_col33[1] <= fa_s4_c33_n15_s;
                    stage5_col33[2] <= stage4_col33[3];
                    stage5_col34[0] <= fa_s4_c33_n15_c;
                    stage5_col34[1] <= fa_s4_c34_n16_s;
                    stage5_col34[2] <= stage4_col34[3];
                    stage5_col35[0] <= fa_s4_c34_n16_c;
                    stage5_col35[1] <= fa_s4_c35_n17_s;
                    stage5_col35[2] <= stage4_col35[3];
                    stage5_col36[0] <= fa_s4_c35_n17_c;
                    stage5_col36[1] <= fa_s4_c36_n18_s;
                    stage5_col36[2] <= stage4_col36[3];
                    stage5_col37[0] <= fa_s4_c36_n18_c;
                    stage5_col37[1] <= fa_s4_c37_n19_s;
                    stage5_col37[2] <= stage4_col37[3];
                    stage5_col38[0] <= fa_s4_c37_n19_c;
                    stage5_col38[1] <= fa_s4_c38_n20_s;
                    stage5_col38[2] <= stage4_col38[3];
                    stage5_col39[0] <= fa_s4_c38_n20_c;
                    stage5_col39[1] <= fa_s4_c39_n21_s;
                    stage5_col39[2] <= stage4_col39[3];
                    stage5_col40[0] <= fa_s4_c39_n21_c;
                    stage5_col40[1] <= fa_s4_c40_n22_s;
                    stage5_col40[2] <= fa_s4_c40_n23_s;
                    stage5_col41[0] <= fa_s4_c40_n22_c;
                    stage5_col41[1] <= fa_s4_c40_n23_c;
                    stage5_col41[2] <= fa_s4_c41_n24_s;
                    stage5_col41[3] <= stage4_col41[3];
                    stage5_col41[4] <= stage4_col41[4];
                    stage5_col42[0] <= fa_s4_c41_n24_c;
                    stage5_col42[1] <= fa_s4_c42_n25_s;
                    stage5_col42[2] <= stage4_col42[3];
                    stage5_col42[3] <= stage4_col42[4];
                    stage5_col43[0] <= fa_s4_c42_n25_c;
                    stage5_col43[1] <= fa_s4_c43_n26_s;
                    stage5_col43[2] <= stage4_col43[3];
                    stage5_col43[3] <= stage4_col43[4];
                    stage5_col44[0] <= fa_s4_c43_n26_c;
                    stage5_col44[1] <= fa_s4_c44_n27_s;
                    stage5_col44[2] <= stage4_col44[3];
                    stage5_col44[3] <= stage4_col44[4];
                    stage5_col45[0] <= fa_s4_c44_n27_c;
                    stage5_col45[1] <= fa_s4_c45_n28_s;
                    stage5_col45[2] <= stage4_col45[3];
                    stage5_col45[3] <= stage4_col45[4];
                    stage5_col46[0] <= fa_s4_c45_n28_c;
                    stage5_col46[1] <= fa_s4_c46_n29_s;
                    stage5_col46[2] <= stage4_col46[3];
                    stage5_col46[3] <= stage4_col46[4];
                    stage5_col47[0] <= fa_s4_c46_n29_c;
                    stage5_col47[1] <= fa_s4_c47_n30_s;
                    stage5_col47[2] <= fa_s4_c47_n31_s;
                    stage5_col47[3] <= stage4_col47[6];
                    stage5_col48[0] <= fa_s4_c47_n30_c;
                    stage5_col48[1] <= fa_s4_c47_n31_c;
                    stage5_col48[2] <= fa_s4_c48_n32_s;
                    stage5_col48[3] <= fa_s4_c48_n33_s;
                    stage5_col49[0] <= fa_s4_c48_n32_c;
                    stage5_col49[1] <= fa_s4_c48_n33_c;
                    stage5_col49[2] <= fa_s4_c49_n34_s;
                    stage5_col49[3] <= fa_s4_c49_n35_s;
                    stage5_col50[0] <= fa_s4_c49_n34_c;
                    stage5_col50[1] <= fa_s4_c49_n35_c;
                    stage5_col50[2] <= fa_s4_c50_n36_s;
                    stage5_col50[3] <= fa_s4_c50_n37_s;
                    stage5_col51[0] <= fa_s4_c50_n36_c;
                    stage5_col51[1] <= fa_s4_c50_n37_c;
                    stage5_col51[2] <= fa_s4_c51_n38_s;
                    stage5_col51[3] <= fa_s4_c51_n39_s;
                    stage5_col52[0] <= fa_s4_c51_n38_c;
                    stage5_col52[1] <= fa_s4_c51_n39_c;
                    stage5_col52[2] <= fa_s4_c52_n40_s;
                    stage5_col52[3] <= fa_s4_c52_n41_s;
                    stage5_col53[0] <= fa_s4_c52_n40_c;
                    stage5_col53[1] <= fa_s4_c52_n41_c;
                    stage5_col53[2] <= fa_s4_c53_n42_s;
                    stage5_col53[3] <= fa_s4_c53_n43_s;
                    stage5_col54[0] <= fa_s4_c53_n42_c;
                    stage5_col54[1] <= fa_s4_c53_n43_c;
                    stage5_col54[2] <= fa_s4_c54_n44_s;
                    stage5_col54[3] <= fa_s4_c54_n45_s;
                    stage5_col55[0] <= fa_s4_c54_n44_c;
                    stage5_col55[1] <= fa_s4_c54_n45_c;
                    stage5_col55[2] <= fa_s4_c55_n46_s;
                    stage5_col55[3] <= fa_s4_c55_n47_s;
                    stage5_col56[0] <= fa_s4_c55_n46_c;
                    stage5_col56[1] <= fa_s4_c55_n47_c;
                    stage5_col56[2] <= fa_s4_c56_n48_s;
                    stage5_col56[3] <= fa_s4_c56_n49_s;
                    stage5_col57[0] <= fa_s4_c56_n48_c;
                    stage5_col57[1] <= fa_s4_c56_n49_c;
                    stage5_col57[2] <= fa_s4_c57_n50_s;
                    stage5_col57[3] <= fa_s4_c57_n51_s;
                    stage5_col58[0] <= fa_s4_c57_n50_c;
                    stage5_col58[1] <= fa_s4_c57_n51_c;
                    stage5_col58[2] <= fa_s4_c58_n52_s;
                    stage5_col58[3] <= fa_s4_c58_n53_s;
                    stage5_col59[0] <= fa_s4_c58_n52_c;
                    stage5_col59[1] <= fa_s4_c58_n53_c;
                    stage5_col59[2] <= fa_s4_c59_n54_s;
                    stage5_col59[3] <= fa_s4_c59_n55_s;
                    stage5_col59[4] <= stage4_col59[6];
                    stage5_col59[5] <= stage4_col59[7];
                    stage5_col60[0] <= fa_s4_c59_n54_c;
                    stage5_col60[1] <= fa_s4_c59_n55_c;
                    stage5_col60[2] <= fa_s4_c60_n56_s;
                    stage5_col60[3] <= fa_s4_c60_n57_s;
                    stage5_col60[4] <= stage4_col60[6];
                    stage5_col61[0] <= fa_s4_c60_n56_c;
                    stage5_col61[1] <= fa_s4_c60_n57_c;
                    stage5_col61[2] <= fa_s4_c61_n58_s;
                    stage5_col61[3] <= fa_s4_c61_n59_s;
                    stage5_col61[4] <= stage4_col61[6];
                    stage5_col62[0] <= fa_s4_c61_n58_c;
                    stage5_col62[1] <= fa_s4_c61_n59_c;
                    stage5_col62[2] <= fa_s4_c62_n60_s;
                    stage5_col62[3] <= fa_s4_c62_n61_s;
                    stage5_col62[4] <= stage4_col62[6];
                    stage5_col63[0] <= fa_s4_c62_n60_c;
                    stage5_col63[1] <= fa_s4_c62_n61_c;
                    stage5_col63[2] <= fa_s4_c63_n62_s;
                    stage5_col63[3] <= fa_s4_c63_n63_s;
                    stage5_col63[4] <= stage4_col63[6];
                    stage5_col64[0] <= fa_s4_c63_n62_c;
                    stage5_col64[1] <= fa_s4_c63_n63_c;
                    stage5_col64[2] <= fa_s4_c64_n64_s;
                    stage5_col64[3] <= fa_s4_c64_n65_s;
                    stage5_col64[4] <= stage4_col64[6];
                    stage5_col64[5] <= stage4_col64[7];
                    stage5_col65[0] <= fa_s4_c64_n64_c;
                    stage5_col65[1] <= fa_s4_c64_n65_c;
                    stage5_col65[2] <= fa_s4_c65_n66_s;
                    stage5_col65[3] <= fa_s4_c65_n67_s;
                    stage5_col65[4] <= stage4_col65[6];
                    stage5_col66[0] <= fa_s4_c65_n66_c;
                    stage5_col66[1] <= fa_s4_c65_n67_c;
                    stage5_col66[2] <= fa_s4_c66_n68_s;
                    stage5_col66[3] <= fa_s4_c66_n69_s;
                    stage5_col66[4] <= stage4_col66[6];
                    stage5_col66[5] <= stage4_col66[7];
                    stage5_col67[0] <= fa_s4_c66_n68_c;
                    stage5_col67[1] <= fa_s4_c66_n69_c;
                    stage5_col67[2] <= fa_s4_c67_n70_s;
                    stage5_col67[3] <= fa_s4_c67_n71_s;
                    stage5_col67[4] <= stage4_col67[6];
                    stage5_col68[0] <= fa_s4_c67_n70_c;
                    stage5_col68[1] <= fa_s4_c67_n71_c;
                    stage5_col68[2] <= fa_s4_c68_n72_s;
                    stage5_col68[3] <= fa_s4_c68_n73_s;
                    stage5_col68[4] <= stage4_col68[6];
                    stage5_col68[5] <= stage4_col68[7];
                    stage5_col69[0] <= fa_s4_c68_n72_c;
                    stage5_col69[1] <= fa_s4_c68_n73_c;
                    stage5_col69[2] <= fa_s4_c69_n74_s;
                    stage5_col69[3] <= fa_s4_c69_n75_s;
                    stage5_col69[4] <= stage4_col69[6];
                    stage5_col70[0] <= fa_s4_c69_n74_c;
                    stage5_col70[1] <= fa_s4_c69_n75_c;
                    stage5_col70[2] <= fa_s4_c70_n76_s;
                    stage5_col70[3] <= fa_s4_c70_n77_s;
                    stage5_col70[4] <= stage4_col70[6];
                    stage5_col70[5] <= stage4_col70[7];
                    stage5_col71[0] <= fa_s4_c70_n76_c;
                    stage5_col71[1] <= fa_s4_c70_n77_c;
                    stage5_col71[2] <= fa_s4_c71_n78_s;
                    stage5_col71[3] <= fa_s4_c71_n79_s;
                    stage5_col71[4] <= stage4_col71[6];
                    stage5_col72[0] <= fa_s4_c71_n78_c;
                    stage5_col72[1] <= fa_s4_c71_n79_c;
                    stage5_col72[2] <= fa_s4_c72_n80_s;
                    stage5_col72[3] <= fa_s4_c72_n81_s;
                    stage5_col72[4] <= stage4_col72[6];
                    stage5_col72[5] <= stage4_col72[7];
                    stage5_col73[0] <= fa_s4_c72_n80_c;
                    stage5_col73[1] <= fa_s4_c72_n81_c;
                    stage5_col73[2] <= fa_s4_c73_n82_s;
                    stage5_col73[3] <= fa_s4_c73_n83_s;
                    stage5_col73[4] <= stage4_col73[6];
                    stage5_col74[0] <= fa_s4_c73_n82_c;
                    stage5_col74[1] <= fa_s4_c73_n83_c;
                    stage5_col74[2] <= fa_s4_c74_n84_s;
                    stage5_col74[3] <= fa_s4_c74_n85_s;
                    stage5_col74[4] <= stage4_col74[6];
                    stage5_col74[5] <= stage4_col74[7];
                    stage5_col75[0] <= fa_s4_c74_n84_c;
                    stage5_col75[1] <= fa_s4_c74_n85_c;
                    stage5_col75[2] <= fa_s4_c75_n86_s;
                    stage5_col75[3] <= fa_s4_c75_n87_s;
                    stage5_col75[4] <= stage4_col75[6];
                    stage5_col76[0] <= fa_s4_c75_n86_c;
                    stage5_col76[1] <= fa_s4_c75_n87_c;
                    stage5_col76[2] <= fa_s4_c76_n88_s;
                    stage5_col76[3] <= fa_s4_c76_n89_s;
                    stage5_col76[4] <= stage4_col76[6];
                    stage5_col76[5] <= stage4_col76[7];
                    stage5_col77[0] <= fa_s4_c76_n88_c;
                    stage5_col77[1] <= fa_s4_c76_n89_c;
                    stage5_col77[2] <= fa_s4_c77_n90_s;
                    stage5_col77[3] <= fa_s4_c77_n91_s;
                    stage5_col77[4] <= stage4_col77[6];
                    stage5_col78[0] <= fa_s4_c77_n90_c;
                    stage5_col78[1] <= fa_s4_c77_n91_c;
                    stage5_col78[2] <= fa_s4_c78_n92_s;
                    stage5_col78[3] <= fa_s4_c78_n93_s;
                    stage5_col78[4] <= stage4_col78[6];
                    stage5_col78[5] <= stage4_col78[7];
                    stage5_col79[0] <= fa_s4_c78_n92_c;
                    stage5_col79[1] <= fa_s4_c78_n93_c;
                    stage5_col79[2] <= fa_s4_c79_n94_s;
                    stage5_col79[3] <= fa_s4_c79_n95_s;
                    stage5_col79[4] <= stage4_col79[6];
                    stage5_col80[0] <= fa_s4_c79_n94_c;
                    stage5_col80[1] <= fa_s4_c79_n95_c;
                    stage5_col80[2] <= fa_s4_c80_n96_s;
                    stage5_col80[3] <= fa_s4_c80_n97_s;
                    stage5_col80[4] <= stage4_col80[6];
                    stage5_col80[5] <= stage4_col80[7];
                    stage5_col81[0] <= fa_s4_c80_n96_c;
                    stage5_col81[1] <= fa_s4_c80_n97_c;
                    stage5_col81[2] <= fa_s4_c81_n98_s;
                    stage5_col81[3] <= fa_s4_c81_n99_s;
                    stage5_col81[4] <= stage4_col81[6];
                    stage5_col82[0] <= fa_s4_c81_n98_c;
                    stage5_col82[1] <= fa_s4_c81_n99_c;
                    stage5_col82[2] <= fa_s4_c82_n100_s;
                    stage5_col82[3] <= fa_s4_c82_n101_s;
                    stage5_col82[4] <= stage4_col82[6];
                    stage5_col82[5] <= stage4_col82[7];
                    stage5_col83[0] <= fa_s4_c82_n100_c;
                    stage5_col83[1] <= fa_s4_c82_n101_c;
                    stage5_col83[2] <= fa_s4_c83_n102_s;
                    stage5_col83[3] <= fa_s4_c83_n103_s;
                    stage5_col83[4] <= stage4_col83[6];
                    stage5_col84[0] <= fa_s4_c83_n102_c;
                    stage5_col84[1] <= fa_s4_c83_n103_c;
                    stage5_col84[2] <= fa_s4_c84_n104_s;
                    stage5_col84[3] <= fa_s4_c84_n105_s;
                    stage5_col84[4] <= stage4_col84[6];
                    stage5_col84[5] <= stage4_col84[7];
                    stage5_col85[0] <= fa_s4_c84_n104_c;
                    stage5_col85[1] <= fa_s4_c84_n105_c;
                    stage5_col85[2] <= fa_s4_c85_n106_s;
                    stage5_col85[3] <= fa_s4_c85_n107_s;
                    stage5_col85[4] <= stage4_col85[6];
                    stage5_col86[0] <= fa_s4_c85_n106_c;
                    stage5_col86[1] <= fa_s4_c85_n107_c;
                    stage5_col86[2] <= fa_s4_c86_n108_s;
                    stage5_col86[3] <= fa_s4_c86_n109_s;
                    stage5_col86[4] <= stage4_col86[6];
                    stage5_col86[5] <= stage4_col86[7];
                    stage5_col87[0] <= fa_s4_c86_n108_c;
                    stage5_col87[1] <= fa_s4_c86_n109_c;
                    stage5_col87[2] <= fa_s4_c87_n110_s;
                    stage5_col87[3] <= fa_s4_c87_n111_s;
                    stage5_col87[4] <= stage4_col87[6];
                    stage5_col88[0] <= fa_s4_c87_n110_c;
                    stage5_col88[1] <= fa_s4_c87_n111_c;
                    stage5_col88[2] <= fa_s4_c88_n112_s;
                    stage5_col88[3] <= fa_s4_c88_n113_s;
                    stage5_col88[4] <= stage4_col88[6];
                    stage5_col88[5] <= stage4_col88[7];
                    stage5_col89[0] <= fa_s4_c88_n112_c;
                    stage5_col89[1] <= fa_s4_c88_n113_c;
                    stage5_col89[2] <= fa_s4_c89_n114_s;
                    stage5_col89[3] <= fa_s4_c89_n115_s;
                    stage5_col89[4] <= stage4_col89[6];
                    stage5_col90[0] <= fa_s4_c89_n114_c;
                    stage5_col90[1] <= fa_s4_c89_n115_c;
                    stage5_col90[2] <= fa_s4_c90_n116_s;
                    stage5_col90[3] <= fa_s4_c90_n117_s;
                    stage5_col90[4] <= stage4_col90[6];
                    stage5_col90[5] <= stage4_col90[7];
                    stage5_col91[0] <= fa_s4_c90_n116_c;
                    stage5_col91[1] <= fa_s4_c90_n117_c;
                    stage5_col91[2] <= fa_s4_c91_n118_s;
                    stage5_col91[3] <= fa_s4_c91_n119_s;
                    stage5_col91[4] <= stage4_col91[6];
                    stage5_col92[0] <= fa_s4_c91_n118_c;
                    stage5_col92[1] <= fa_s4_c91_n119_c;
                    stage5_col92[2] <= fa_s4_c92_n120_s;
                    stage5_col92[3] <= fa_s4_c92_n121_s;
                    stage5_col92[4] <= stage4_col92[6];
                    stage5_col92[5] <= stage4_col92[7];
                    stage5_col93[0] <= fa_s4_c92_n120_c;
                    stage5_col93[1] <= fa_s4_c92_n121_c;
                    stage5_col93[2] <= fa_s4_c93_n122_s;
                    stage5_col93[3] <= fa_s4_c93_n123_s;
                    stage5_col93[4] <= stage4_col93[6];
                    stage5_col94[0] <= fa_s4_c93_n122_c;
                    stage5_col94[1] <= fa_s4_c93_n123_c;
                    stage5_col94[2] <= fa_s4_c94_n124_s;
                    stage5_col94[3] <= fa_s4_c94_n125_s;
                    stage5_col94[4] <= stage4_col94[6];
                    stage5_col94[5] <= stage4_col94[7];
                    stage5_col95[0] <= fa_s4_c94_n124_c;
                    stage5_col95[1] <= fa_s4_c94_n125_c;
                    stage5_col95[2] <= fa_s4_c95_n126_s;
                    stage5_col95[3] <= fa_s4_c95_n127_s;
                    stage5_col95[4] <= stage4_col95[6];
                    stage5_col96[0] <= fa_s4_c95_n126_c;
                    stage5_col96[1] <= fa_s4_c95_n127_c;
                    stage5_col96[2] <= fa_s4_c96_n128_s;
                    stage5_col96[3] <= fa_s4_c96_n129_s;
                    stage5_col96[4] <= stage4_col96[6];
                    stage5_col96[5] <= stage4_col96[7];
                    stage5_col97[0] <= fa_s4_c96_n128_c;
                    stage5_col97[1] <= fa_s4_c96_n129_c;
                    stage5_col97[2] <= fa_s4_c97_n130_s;
                    stage5_col97[3] <= fa_s4_c97_n131_s;
                    stage5_col97[4] <= stage4_col97[6];
                    stage5_col98[0] <= fa_s4_c97_n130_c;
                    stage5_col98[1] <= fa_s4_c97_n131_c;
                    stage5_col98[2] <= fa_s4_c98_n132_s;
                    stage5_col98[3] <= fa_s4_c98_n133_s;
                    stage5_col98[4] <= stage4_col98[6];
                    stage5_col98[5] <= stage4_col98[7];
                    stage5_col99[0] <= fa_s4_c98_n132_c;
                    stage5_col99[1] <= fa_s4_c98_n133_c;
                    stage5_col99[2] <= fa_s4_c99_n134_s;
                    stage5_col99[3] <= fa_s4_c99_n135_s;
                    stage5_col99[4] <= stage4_col99[6];
                    stage5_col100[0] <= fa_s4_c99_n134_c;
                    stage5_col100[1] <= fa_s4_c99_n135_c;
                    stage5_col100[2] <= fa_s4_c100_n136_s;
                    stage5_col100[3] <= fa_s4_c100_n137_s;
                    stage5_col100[4] <= stage4_col100[6];
                    stage5_col100[5] <= stage4_col100[7];
                    stage5_col101[0] <= fa_s4_c100_n136_c;
                    stage5_col101[1] <= fa_s4_c100_n137_c;
                    stage5_col101[2] <= fa_s4_c101_n138_s;
                    stage5_col101[3] <= fa_s4_c101_n139_s;
                    stage5_col101[4] <= stage4_col101[6];
                    stage5_col102[0] <= fa_s4_c101_n138_c;
                    stage5_col102[1] <= fa_s4_c101_n139_c;
                    stage5_col102[2] <= fa_s4_c102_n140_s;
                    stage5_col102[3] <= fa_s4_c102_n141_s;
                    stage5_col102[4] <= stage4_col102[6];
                    stage5_col102[5] <= stage4_col102[7];
                    stage5_col103[0] <= fa_s4_c102_n140_c;
                    stage5_col103[1] <= fa_s4_c102_n141_c;
                    stage5_col103[2] <= fa_s4_c103_n142_s;
                    stage5_col103[3] <= fa_s4_c103_n143_s;
                    stage5_col103[4] <= stage4_col103[6];
                    stage5_col104[0] <= fa_s4_c103_n142_c;
                    stage5_col104[1] <= fa_s4_c103_n143_c;
                    stage5_col104[2] <= fa_s4_c104_n144_s;
                    stage5_col104[3] <= fa_s4_c104_n145_s;
                    stage5_col104[4] <= stage4_col104[6];
                    stage5_col104[5] <= stage4_col104[7];
                    stage5_col105[0] <= fa_s4_c104_n144_c;
                    stage5_col105[1] <= fa_s4_c104_n145_c;
                    stage5_col105[2] <= fa_s4_c105_n146_s;
                    stage5_col105[3] <= fa_s4_c105_n147_s;
                    stage5_col105[4] <= stage4_col105[6];
                    stage5_col106[0] <= fa_s4_c105_n146_c;
                    stage5_col106[1] <= fa_s4_c105_n147_c;
                    stage5_col106[2] <= fa_s4_c106_n148_s;
                    stage5_col106[3] <= fa_s4_c106_n149_s;
                    stage5_col106[4] <= stage4_col106[6];
                    stage5_col106[5] <= stage4_col106[7];
                    stage5_col107[0] <= fa_s4_c106_n148_c;
                    stage5_col107[1] <= fa_s4_c106_n149_c;
                    stage5_col107[2] <= fa_s4_c107_n150_s;
                    stage5_col107[3] <= fa_s4_c107_n151_s;
                    stage5_col107[4] <= stage4_col107[6];
                    stage5_col108[0] <= fa_s4_c107_n150_c;
                    stage5_col108[1] <= fa_s4_c107_n151_c;
                    stage5_col108[2] <= fa_s4_c108_n152_s;
                    stage5_col108[3] <= fa_s4_c108_n153_s;
                    stage5_col108[4] <= stage4_col108[6];
                    stage5_col108[5] <= stage4_col108[7];
                    stage5_col109[0] <= fa_s4_c108_n152_c;
                    stage5_col109[1] <= fa_s4_c108_n153_c;
                    stage5_col109[2] <= fa_s4_c109_n154_s;
                    stage5_col109[3] <= fa_s4_c109_n155_s;
                    stage5_col109[4] <= stage4_col109[6];
                    stage5_col110[0] <= fa_s4_c109_n154_c;
                    stage5_col110[1] <= fa_s4_c109_n155_c;
                    stage5_col110[2] <= fa_s4_c110_n156_s;
                    stage5_col110[3] <= fa_s4_c110_n157_s;
                    stage5_col110[4] <= stage4_col110[6];
                    stage5_col110[5] <= stage4_col110[7];
                    stage5_col111[0] <= fa_s4_c110_n156_c;
                    stage5_col111[1] <= fa_s4_c110_n157_c;
                    stage5_col111[2] <= fa_s4_c111_n158_s;
                    stage5_col111[3] <= fa_s4_c111_n159_s;
                    stage5_col111[4] <= stage4_col111[6];
                    stage5_col112[0] <= fa_s4_c111_n158_c;
                    stage5_col112[1] <= fa_s4_c111_n159_c;
                    stage5_col112[2] <= fa_s4_c112_n160_s;
                    stage5_col112[3] <= fa_s4_c112_n161_s;
                    stage5_col112[4] <= stage4_col112[6];
                    stage5_col112[5] <= stage4_col112[7];
                    stage5_col113[0] <= fa_s4_c112_n160_c;
                    stage5_col113[1] <= fa_s4_c112_n161_c;
                    stage5_col113[2] <= fa_s4_c113_n162_s;
                    stage5_col113[3] <= fa_s4_c113_n163_s;
                    stage5_col113[4] <= stage4_col113[6];
                    stage5_col114[0] <= fa_s4_c113_n162_c;
                    stage5_col114[1] <= fa_s4_c113_n163_c;
                    stage5_col114[2] <= fa_s4_c114_n164_s;
                    stage5_col114[3] <= fa_s4_c114_n165_s;
                    stage5_col114[4] <= stage4_col114[6];
                    stage5_col114[5] <= stage4_col114[7];
                    stage5_col115[0] <= fa_s4_c114_n164_c;
                    stage5_col115[1] <= fa_s4_c114_n165_c;
                    stage5_col115[2] <= fa_s4_c115_n166_s;
                    stage5_col115[3] <= fa_s4_c115_n167_s;
                    stage5_col115[4] <= stage4_col115[6];
                    stage5_col116[0] <= fa_s4_c115_n166_c;
                    stage5_col116[1] <= fa_s4_c115_n167_c;
                    stage5_col116[2] <= fa_s4_c116_n168_s;
                    stage5_col116[3] <= fa_s4_c116_n169_s;
                    stage5_col116[4] <= stage4_col116[6];
                    stage5_col116[5] <= stage4_col116[7];
                    stage5_col117[0] <= fa_s4_c116_n168_c;
                    stage5_col117[1] <= fa_s4_c116_n169_c;
                    stage5_col117[2] <= fa_s4_c117_n170_s;
                    stage5_col117[3] <= fa_s4_c117_n171_s;
                    stage5_col117[4] <= stage4_col117[6];
                    stage5_col118[0] <= fa_s4_c117_n170_c;
                    stage5_col118[1] <= fa_s4_c117_n171_c;
                    stage5_col118[2] <= fa_s4_c118_n172_s;
                    stage5_col118[3] <= fa_s4_c118_n173_s;
                    stage5_col118[4] <= stage4_col118[6];
                    stage5_col118[5] <= stage4_col118[7];
                    stage5_col119[0] <= fa_s4_c118_n172_c;
                    stage5_col119[1] <= fa_s4_c118_n173_c;
                    stage5_col119[2] <= fa_s4_c119_n174_s;
                    stage5_col119[3] <= fa_s4_c119_n175_s;
                    stage5_col119[4] <= stage4_col119[6];
                    stage5_col120[0] <= fa_s4_c119_n174_c;
                    stage5_col120[1] <= fa_s4_c119_n175_c;
                    stage5_col120[2] <= fa_s4_c120_n176_s;
                    stage5_col120[3] <= fa_s4_c120_n177_s;
                    stage5_col120[4] <= stage4_col120[6];
                    stage5_col120[5] <= stage4_col120[7];
                    stage5_col121[0] <= fa_s4_c120_n176_c;
                    stage5_col121[1] <= fa_s4_c120_n177_c;
                    stage5_col121[2] <= fa_s4_c121_n178_s;
                    stage5_col121[3] <= fa_s4_c121_n179_s;
                    stage5_col121[4] <= stage4_col121[6];
                    stage5_col122[0] <= fa_s4_c121_n178_c;
                    stage5_col122[1] <= fa_s4_c121_n179_c;
                    stage5_col122[2] <= fa_s4_c122_n180_s;
                    stage5_col122[3] <= fa_s4_c122_n181_s;
                    stage5_col122[4] <= stage4_col122[6];
                    stage5_col122[5] <= stage4_col122[7];
                    stage5_col123[0] <= fa_s4_c122_n180_c;
                    stage5_col123[1] <= fa_s4_c122_n181_c;
                    stage5_col123[2] <= fa_s4_c123_n182_s;
                    stage5_col123[3] <= fa_s4_c123_n183_s;
                    stage5_col123[4] <= stage4_col123[6];
                    stage5_col124[0] <= fa_s4_c123_n182_c;
                    stage5_col124[1] <= fa_s4_c123_n183_c;
                    stage5_col124[2] <= fa_s4_c124_n184_s;
                    stage5_col124[3] <= fa_s4_c124_n185_s;
                    stage5_col124[4] <= stage4_col124[6];
                    stage5_col124[5] <= stage4_col124[7];
                    stage5_col125[0] <= fa_s4_c124_n184_c;
                    stage5_col125[1] <= fa_s4_c124_n185_c;
                    stage5_col125[2] <= fa_s4_c125_n186_s;
                    stage5_col125[3] <= fa_s4_c125_n187_s;
                    stage5_col125[4] <= stage4_col125[6];
                    stage5_col126[0] <= fa_s4_c125_n186_c;
                    stage5_col126[1] <= fa_s4_c125_n187_c;
                    stage5_col126[2] <= fa_s4_c126_n188_s;
                    stage5_col126[3] <= fa_s4_c126_n189_s;
                    stage5_col126[4] <= stage4_col126[6];
                    stage5_col126[5] <= stage4_col126[7];
                    stage5_col127[0] <= fa_s4_c126_n188_c;
                    stage5_col127[1] <= fa_s4_c126_n189_c;
                    stage5_col127[2] <= stage4_col127[0];
                    stage5_col127[3] <= stage4_col127[1];
                    stage5_col127[4] <= stage4_col127[2];
                    stage5_col127[5] <= stage4_col127[3];
                    stage5_col127[6] <= stage4_col127[4];
                    stage5_col127[7] <= stage4_col127[5];
                    stage5_col127[8] <= stage4_col127[6];
                    stage5_col127[9] <= stage4_col127[7];
                    stage5_col127[10] <= stage4_col127[8];
                    stage5_col127[11] <= stage4_col127[9];
                    stage5_col127[12] <= stage4_col127[10];
                    stage5_col127[13] <= stage4_col127[11];
                    stage5_col127[14] <= stage4_col127[12];
                    stage5_col127[15] <= stage4_col127[13];
                    stage5_col127[16] <= stage4_col127[14];
                    stage5_col127[17] <= stage4_col127[15];
                    stage5_col127[18] <= stage4_col127[16];
                    stage5_col127[19] <= stage4_col127[17];
                    stage5_col127[20] <= stage4_col127[18];
                    stage5_col127[21] <= stage4_col127[19];
                    stage5_col127[22] <= stage4_col127[20];
                    stage5_col127[23] <= stage4_col127[21];
                    stage5_col127[24] <= stage4_col127[22];
                    stage5_col127[25] <= stage4_col127[23];
                    stage5_col127[26] <= stage4_col127[24];
                    stage5_col127[27] <= stage4_col127[25];
                    stage5_col127[28] <= stage4_col127[25];
                    stage5_col127[29] <= stage4_col127[25];
                    stage5_col127[30] <= stage4_col127[25];
                    stage5_col127[31] <= stage4_col127[25];
                    stage5_col127[32] <= stage4_col127[25];
                    stage5_col127[33] <= stage4_col127[25];
                    stage5_col127[34] <= stage4_col127[25];
                    stage5_col127[35] <= stage4_col127[25];
                    stage5_col127[36] <= stage4_col127[25];
                    stage5_col127[37] <= stage4_col127[25];
                    stage5_col127[38] <= stage4_col127[25];
                    stage5_col127[39] <= stage4_col127[25];
                    stage5_col127[40] <= stage4_col127[25];
                    stage5_col127[41] <= stage4_col127[25];
                    stage5_col127[42] <= stage4_col127[25];
                    stage5_col127[43] <= stage4_col127[25];
                    stage5_col127[44] <= stage4_col127[25];
                    stage5_col127[45] <= stage4_col127[25];
                    stage5_col127[46] <= stage4_col127[25];
                    stage5_col127[47] <= stage4_col127[25];
                    stage5_col127[48] <= stage4_col127[25];
                    stage5_col127[49] <= stage4_col127[25];
                    stage5_col127[50] <= stage4_col127[25];
                    stage5_col127[51] <= stage4_col127[25];
                    stage5_col127[52] <= stage4_col127[25];
                    stage5_col127[53] <= stage4_col127[25];
                    stage5_col127[54] <= stage4_col127[25];
                    stage5_col127[55] <= stage4_col127[25];
                    stage5_col127[56] <= stage4_col127[25];
                    stage5_col127[57] <= stage4_col127[25];
                    stage5_col127[58] <= stage4_col127[25];
                end
            end
        end else begin : gen_stage5_no_pipe
            // Combinational assignment
            always_comb begin
                stage5_col0[0] = stage4_col0[0];
                stage5_col1[0] = stage4_col1[0];
                stage5_col2[0] = stage4_col2[0];
                stage5_col3[0] = stage4_col3[0];
                stage5_col4[0] = ha_s4_c4_n0_s;
                stage5_col5[0] = ha_s4_c4_n0_c;
                stage5_col5[1] = stage4_col5[0];
                stage5_col6[0] = fa_s4_c6_n0_s;
                stage5_col7[0] = fa_s4_c6_n0_c;
                stage5_col7[1] = stage4_col7[0];
                stage5_col7[2] = stage4_col7[1];
                stage5_col8[0] = stage4_col8[0];
                stage5_col8[1] = stage4_col8[1];
                stage5_col9[0] = stage4_col9[0];
                stage5_col9[1] = stage4_col9[1];
                stage5_col10[0] = stage4_col10[0];
                stage5_col10[1] = stage4_col10[1];
                stage5_col11[0] = stage4_col11[0];
                stage5_col11[1] = stage4_col11[1];
                stage5_col12[0] = stage4_col12[0];
                stage5_col12[1] = stage4_col12[1];
                stage5_col13[0] = stage4_col13[0];
                stage5_col13[1] = stage4_col13[1];
                stage5_col14[0] = stage4_col14[0];
                stage5_col14[1] = stage4_col14[1];
                stage5_col15[0] = stage4_col15[0];
                stage5_col15[1] = stage4_col15[1];
                stage5_col16[0] = stage4_col16[0];
                stage5_col16[1] = stage4_col16[1];
                stage5_col17[0] = stage4_col17[0];
                stage5_col17[1] = stage4_col17[1];
                stage5_col18[0] = stage4_col18[0];
                stage5_col18[1] = stage4_col18[1];
                stage5_col19[0] = fa_s4_c19_n1_s;
                stage5_col19[1] = stage4_col19[3];
                stage5_col20[0] = fa_s4_c19_n1_c;
                stage5_col20[1] = fa_s4_c20_n2_s;
                stage5_col21[0] = fa_s4_c20_n2_c;
                stage5_col21[1] = fa_s4_c21_n3_s;
                stage5_col22[0] = fa_s4_c21_n3_c;
                stage5_col22[1] = fa_s4_c22_n4_s;
                stage5_col23[0] = fa_s4_c22_n4_c;
                stage5_col23[1] = fa_s4_c23_n5_s;
                stage5_col24[0] = fa_s4_c23_n5_c;
                stage5_col24[1] = fa_s4_c24_n6_s;
                stage5_col25[0] = fa_s4_c24_n6_c;
                stage5_col25[1] = fa_s4_c25_n7_s;
                stage5_col26[0] = fa_s4_c25_n7_c;
                stage5_col26[1] = fa_s4_c26_n8_s;
                stage5_col27[0] = fa_s4_c26_n8_c;
                stage5_col27[1] = fa_s4_c27_n9_s;
                stage5_col28[0] = fa_s4_c27_n9_c;
                stage5_col28[1] = fa_s4_c28_n10_s;
                stage5_col28[2] = stage4_col28[3];
                stage5_col28[3] = stage4_col28[4];
                stage5_col29[0] = fa_s4_c28_n10_c;
                stage5_col29[1] = fa_s4_c29_n11_s;
                stage5_col29[2] = stage4_col29[3];
                stage5_col30[0] = fa_s4_c29_n11_c;
                stage5_col30[1] = fa_s4_c30_n12_s;
                stage5_col30[2] = stage4_col30[3];
                stage5_col31[0] = fa_s4_c30_n12_c;
                stage5_col31[1] = fa_s4_c31_n13_s;
                stage5_col31[2] = stage4_col31[3];
                stage5_col32[0] = fa_s4_c31_n13_c;
                stage5_col32[1] = fa_s4_c32_n14_s;
                stage5_col32[2] = stage4_col32[3];
                stage5_col33[0] = fa_s4_c32_n14_c;
                stage5_col33[1] = fa_s4_c33_n15_s;
                stage5_col33[2] = stage4_col33[3];
                stage5_col34[0] = fa_s4_c33_n15_c;
                stage5_col34[1] = fa_s4_c34_n16_s;
                stage5_col34[2] = stage4_col34[3];
                stage5_col35[0] = fa_s4_c34_n16_c;
                stage5_col35[1] = fa_s4_c35_n17_s;
                stage5_col35[2] = stage4_col35[3];
                stage5_col36[0] = fa_s4_c35_n17_c;
                stage5_col36[1] = fa_s4_c36_n18_s;
                stage5_col36[2] = stage4_col36[3];
                stage5_col37[0] = fa_s4_c36_n18_c;
                stage5_col37[1] = fa_s4_c37_n19_s;
                stage5_col37[2] = stage4_col37[3];
                stage5_col38[0] = fa_s4_c37_n19_c;
                stage5_col38[1] = fa_s4_c38_n20_s;
                stage5_col38[2] = stage4_col38[3];
                stage5_col39[0] = fa_s4_c38_n20_c;
                stage5_col39[1] = fa_s4_c39_n21_s;
                stage5_col39[2] = stage4_col39[3];
                stage5_col40[0] = fa_s4_c39_n21_c;
                stage5_col40[1] = fa_s4_c40_n22_s;
                stage5_col40[2] = fa_s4_c40_n23_s;
                stage5_col41[0] = fa_s4_c40_n22_c;
                stage5_col41[1] = fa_s4_c40_n23_c;
                stage5_col41[2] = fa_s4_c41_n24_s;
                stage5_col41[3] = stage4_col41[3];
                stage5_col41[4] = stage4_col41[4];
                stage5_col42[0] = fa_s4_c41_n24_c;
                stage5_col42[1] = fa_s4_c42_n25_s;
                stage5_col42[2] = stage4_col42[3];
                stage5_col42[3] = stage4_col42[4];
                stage5_col43[0] = fa_s4_c42_n25_c;
                stage5_col43[1] = fa_s4_c43_n26_s;
                stage5_col43[2] = stage4_col43[3];
                stage5_col43[3] = stage4_col43[4];
                stage5_col44[0] = fa_s4_c43_n26_c;
                stage5_col44[1] = fa_s4_c44_n27_s;
                stage5_col44[2] = stage4_col44[3];
                stage5_col44[3] = stage4_col44[4];
                stage5_col45[0] = fa_s4_c44_n27_c;
                stage5_col45[1] = fa_s4_c45_n28_s;
                stage5_col45[2] = stage4_col45[3];
                stage5_col45[3] = stage4_col45[4];
                stage5_col46[0] = fa_s4_c45_n28_c;
                stage5_col46[1] = fa_s4_c46_n29_s;
                stage5_col46[2] = stage4_col46[3];
                stage5_col46[3] = stage4_col46[4];
                stage5_col47[0] = fa_s4_c46_n29_c;
                stage5_col47[1] = fa_s4_c47_n30_s;
                stage5_col47[2] = fa_s4_c47_n31_s;
                stage5_col47[3] = stage4_col47[6];
                stage5_col48[0] = fa_s4_c47_n30_c;
                stage5_col48[1] = fa_s4_c47_n31_c;
                stage5_col48[2] = fa_s4_c48_n32_s;
                stage5_col48[3] = fa_s4_c48_n33_s;
                stage5_col49[0] = fa_s4_c48_n32_c;
                stage5_col49[1] = fa_s4_c48_n33_c;
                stage5_col49[2] = fa_s4_c49_n34_s;
                stage5_col49[3] = fa_s4_c49_n35_s;
                stage5_col50[0] = fa_s4_c49_n34_c;
                stage5_col50[1] = fa_s4_c49_n35_c;
                stage5_col50[2] = fa_s4_c50_n36_s;
                stage5_col50[3] = fa_s4_c50_n37_s;
                stage5_col51[0] = fa_s4_c50_n36_c;
                stage5_col51[1] = fa_s4_c50_n37_c;
                stage5_col51[2] = fa_s4_c51_n38_s;
                stage5_col51[3] = fa_s4_c51_n39_s;
                stage5_col52[0] = fa_s4_c51_n38_c;
                stage5_col52[1] = fa_s4_c51_n39_c;
                stage5_col52[2] = fa_s4_c52_n40_s;
                stage5_col52[3] = fa_s4_c52_n41_s;
                stage5_col53[0] = fa_s4_c52_n40_c;
                stage5_col53[1] = fa_s4_c52_n41_c;
                stage5_col53[2] = fa_s4_c53_n42_s;
                stage5_col53[3] = fa_s4_c53_n43_s;
                stage5_col54[0] = fa_s4_c53_n42_c;
                stage5_col54[1] = fa_s4_c53_n43_c;
                stage5_col54[2] = fa_s4_c54_n44_s;
                stage5_col54[3] = fa_s4_c54_n45_s;
                stage5_col55[0] = fa_s4_c54_n44_c;
                stage5_col55[1] = fa_s4_c54_n45_c;
                stage5_col55[2] = fa_s4_c55_n46_s;
                stage5_col55[3] = fa_s4_c55_n47_s;
                stage5_col56[0] = fa_s4_c55_n46_c;
                stage5_col56[1] = fa_s4_c55_n47_c;
                stage5_col56[2] = fa_s4_c56_n48_s;
                stage5_col56[3] = fa_s4_c56_n49_s;
                stage5_col57[0] = fa_s4_c56_n48_c;
                stage5_col57[1] = fa_s4_c56_n49_c;
                stage5_col57[2] = fa_s4_c57_n50_s;
                stage5_col57[3] = fa_s4_c57_n51_s;
                stage5_col58[0] = fa_s4_c57_n50_c;
                stage5_col58[1] = fa_s4_c57_n51_c;
                stage5_col58[2] = fa_s4_c58_n52_s;
                stage5_col58[3] = fa_s4_c58_n53_s;
                stage5_col59[0] = fa_s4_c58_n52_c;
                stage5_col59[1] = fa_s4_c58_n53_c;
                stage5_col59[2] = fa_s4_c59_n54_s;
                stage5_col59[3] = fa_s4_c59_n55_s;
                stage5_col59[4] = stage4_col59[6];
                stage5_col59[5] = stage4_col59[7];
                stage5_col60[0] = fa_s4_c59_n54_c;
                stage5_col60[1] = fa_s4_c59_n55_c;
                stage5_col60[2] = fa_s4_c60_n56_s;
                stage5_col60[3] = fa_s4_c60_n57_s;
                stage5_col60[4] = stage4_col60[6];
                stage5_col61[0] = fa_s4_c60_n56_c;
                stage5_col61[1] = fa_s4_c60_n57_c;
                stage5_col61[2] = fa_s4_c61_n58_s;
                stage5_col61[3] = fa_s4_c61_n59_s;
                stage5_col61[4] = stage4_col61[6];
                stage5_col62[0] = fa_s4_c61_n58_c;
                stage5_col62[1] = fa_s4_c61_n59_c;
                stage5_col62[2] = fa_s4_c62_n60_s;
                stage5_col62[3] = fa_s4_c62_n61_s;
                stage5_col62[4] = stage4_col62[6];
                stage5_col63[0] = fa_s4_c62_n60_c;
                stage5_col63[1] = fa_s4_c62_n61_c;
                stage5_col63[2] = fa_s4_c63_n62_s;
                stage5_col63[3] = fa_s4_c63_n63_s;
                stage5_col63[4] = stage4_col63[6];
                stage5_col64[0] = fa_s4_c63_n62_c;
                stage5_col64[1] = fa_s4_c63_n63_c;
                stage5_col64[2] = fa_s4_c64_n64_s;
                stage5_col64[3] = fa_s4_c64_n65_s;
                stage5_col64[4] = stage4_col64[6];
                stage5_col64[5] = stage4_col64[7];
                stage5_col65[0] = fa_s4_c64_n64_c;
                stage5_col65[1] = fa_s4_c64_n65_c;
                stage5_col65[2] = fa_s4_c65_n66_s;
                stage5_col65[3] = fa_s4_c65_n67_s;
                stage5_col65[4] = stage4_col65[6];
                stage5_col66[0] = fa_s4_c65_n66_c;
                stage5_col66[1] = fa_s4_c65_n67_c;
                stage5_col66[2] = fa_s4_c66_n68_s;
                stage5_col66[3] = fa_s4_c66_n69_s;
                stage5_col66[4] = stage4_col66[6];
                stage5_col66[5] = stage4_col66[7];
                stage5_col67[0] = fa_s4_c66_n68_c;
                stage5_col67[1] = fa_s4_c66_n69_c;
                stage5_col67[2] = fa_s4_c67_n70_s;
                stage5_col67[3] = fa_s4_c67_n71_s;
                stage5_col67[4] = stage4_col67[6];
                stage5_col68[0] = fa_s4_c67_n70_c;
                stage5_col68[1] = fa_s4_c67_n71_c;
                stage5_col68[2] = fa_s4_c68_n72_s;
                stage5_col68[3] = fa_s4_c68_n73_s;
                stage5_col68[4] = stage4_col68[6];
                stage5_col68[5] = stage4_col68[7];
                stage5_col69[0] = fa_s4_c68_n72_c;
                stage5_col69[1] = fa_s4_c68_n73_c;
                stage5_col69[2] = fa_s4_c69_n74_s;
                stage5_col69[3] = fa_s4_c69_n75_s;
                stage5_col69[4] = stage4_col69[6];
                stage5_col70[0] = fa_s4_c69_n74_c;
                stage5_col70[1] = fa_s4_c69_n75_c;
                stage5_col70[2] = fa_s4_c70_n76_s;
                stage5_col70[3] = fa_s4_c70_n77_s;
                stage5_col70[4] = stage4_col70[6];
                stage5_col70[5] = stage4_col70[7];
                stage5_col71[0] = fa_s4_c70_n76_c;
                stage5_col71[1] = fa_s4_c70_n77_c;
                stage5_col71[2] = fa_s4_c71_n78_s;
                stage5_col71[3] = fa_s4_c71_n79_s;
                stage5_col71[4] = stage4_col71[6];
                stage5_col72[0] = fa_s4_c71_n78_c;
                stage5_col72[1] = fa_s4_c71_n79_c;
                stage5_col72[2] = fa_s4_c72_n80_s;
                stage5_col72[3] = fa_s4_c72_n81_s;
                stage5_col72[4] = stage4_col72[6];
                stage5_col72[5] = stage4_col72[7];
                stage5_col73[0] = fa_s4_c72_n80_c;
                stage5_col73[1] = fa_s4_c72_n81_c;
                stage5_col73[2] = fa_s4_c73_n82_s;
                stage5_col73[3] = fa_s4_c73_n83_s;
                stage5_col73[4] = stage4_col73[6];
                stage5_col74[0] = fa_s4_c73_n82_c;
                stage5_col74[1] = fa_s4_c73_n83_c;
                stage5_col74[2] = fa_s4_c74_n84_s;
                stage5_col74[3] = fa_s4_c74_n85_s;
                stage5_col74[4] = stage4_col74[6];
                stage5_col74[5] = stage4_col74[7];
                stage5_col75[0] = fa_s4_c74_n84_c;
                stage5_col75[1] = fa_s4_c74_n85_c;
                stage5_col75[2] = fa_s4_c75_n86_s;
                stage5_col75[3] = fa_s4_c75_n87_s;
                stage5_col75[4] = stage4_col75[6];
                stage5_col76[0] = fa_s4_c75_n86_c;
                stage5_col76[1] = fa_s4_c75_n87_c;
                stage5_col76[2] = fa_s4_c76_n88_s;
                stage5_col76[3] = fa_s4_c76_n89_s;
                stage5_col76[4] = stage4_col76[6];
                stage5_col76[5] = stage4_col76[7];
                stage5_col77[0] = fa_s4_c76_n88_c;
                stage5_col77[1] = fa_s4_c76_n89_c;
                stage5_col77[2] = fa_s4_c77_n90_s;
                stage5_col77[3] = fa_s4_c77_n91_s;
                stage5_col77[4] = stage4_col77[6];
                stage5_col78[0] = fa_s4_c77_n90_c;
                stage5_col78[1] = fa_s4_c77_n91_c;
                stage5_col78[2] = fa_s4_c78_n92_s;
                stage5_col78[3] = fa_s4_c78_n93_s;
                stage5_col78[4] = stage4_col78[6];
                stage5_col78[5] = stage4_col78[7];
                stage5_col79[0] = fa_s4_c78_n92_c;
                stage5_col79[1] = fa_s4_c78_n93_c;
                stage5_col79[2] = fa_s4_c79_n94_s;
                stage5_col79[3] = fa_s4_c79_n95_s;
                stage5_col79[4] = stage4_col79[6];
                stage5_col80[0] = fa_s4_c79_n94_c;
                stage5_col80[1] = fa_s4_c79_n95_c;
                stage5_col80[2] = fa_s4_c80_n96_s;
                stage5_col80[3] = fa_s4_c80_n97_s;
                stage5_col80[4] = stage4_col80[6];
                stage5_col80[5] = stage4_col80[7];
                stage5_col81[0] = fa_s4_c80_n96_c;
                stage5_col81[1] = fa_s4_c80_n97_c;
                stage5_col81[2] = fa_s4_c81_n98_s;
                stage5_col81[3] = fa_s4_c81_n99_s;
                stage5_col81[4] = stage4_col81[6];
                stage5_col82[0] = fa_s4_c81_n98_c;
                stage5_col82[1] = fa_s4_c81_n99_c;
                stage5_col82[2] = fa_s4_c82_n100_s;
                stage5_col82[3] = fa_s4_c82_n101_s;
                stage5_col82[4] = stage4_col82[6];
                stage5_col82[5] = stage4_col82[7];
                stage5_col83[0] = fa_s4_c82_n100_c;
                stage5_col83[1] = fa_s4_c82_n101_c;
                stage5_col83[2] = fa_s4_c83_n102_s;
                stage5_col83[3] = fa_s4_c83_n103_s;
                stage5_col83[4] = stage4_col83[6];
                stage5_col84[0] = fa_s4_c83_n102_c;
                stage5_col84[1] = fa_s4_c83_n103_c;
                stage5_col84[2] = fa_s4_c84_n104_s;
                stage5_col84[3] = fa_s4_c84_n105_s;
                stage5_col84[4] = stage4_col84[6];
                stage5_col84[5] = stage4_col84[7];
                stage5_col85[0] = fa_s4_c84_n104_c;
                stage5_col85[1] = fa_s4_c84_n105_c;
                stage5_col85[2] = fa_s4_c85_n106_s;
                stage5_col85[3] = fa_s4_c85_n107_s;
                stage5_col85[4] = stage4_col85[6];
                stage5_col86[0] = fa_s4_c85_n106_c;
                stage5_col86[1] = fa_s4_c85_n107_c;
                stage5_col86[2] = fa_s4_c86_n108_s;
                stage5_col86[3] = fa_s4_c86_n109_s;
                stage5_col86[4] = stage4_col86[6];
                stage5_col86[5] = stage4_col86[7];
                stage5_col87[0] = fa_s4_c86_n108_c;
                stage5_col87[1] = fa_s4_c86_n109_c;
                stage5_col87[2] = fa_s4_c87_n110_s;
                stage5_col87[3] = fa_s4_c87_n111_s;
                stage5_col87[4] = stage4_col87[6];
                stage5_col88[0] = fa_s4_c87_n110_c;
                stage5_col88[1] = fa_s4_c87_n111_c;
                stage5_col88[2] = fa_s4_c88_n112_s;
                stage5_col88[3] = fa_s4_c88_n113_s;
                stage5_col88[4] = stage4_col88[6];
                stage5_col88[5] = stage4_col88[7];
                stage5_col89[0] = fa_s4_c88_n112_c;
                stage5_col89[1] = fa_s4_c88_n113_c;
                stage5_col89[2] = fa_s4_c89_n114_s;
                stage5_col89[3] = fa_s4_c89_n115_s;
                stage5_col89[4] = stage4_col89[6];
                stage5_col90[0] = fa_s4_c89_n114_c;
                stage5_col90[1] = fa_s4_c89_n115_c;
                stage5_col90[2] = fa_s4_c90_n116_s;
                stage5_col90[3] = fa_s4_c90_n117_s;
                stage5_col90[4] = stage4_col90[6];
                stage5_col90[5] = stage4_col90[7];
                stage5_col91[0] = fa_s4_c90_n116_c;
                stage5_col91[1] = fa_s4_c90_n117_c;
                stage5_col91[2] = fa_s4_c91_n118_s;
                stage5_col91[3] = fa_s4_c91_n119_s;
                stage5_col91[4] = stage4_col91[6];
                stage5_col92[0] = fa_s4_c91_n118_c;
                stage5_col92[1] = fa_s4_c91_n119_c;
                stage5_col92[2] = fa_s4_c92_n120_s;
                stage5_col92[3] = fa_s4_c92_n121_s;
                stage5_col92[4] = stage4_col92[6];
                stage5_col92[5] = stage4_col92[7];
                stage5_col93[0] = fa_s4_c92_n120_c;
                stage5_col93[1] = fa_s4_c92_n121_c;
                stage5_col93[2] = fa_s4_c93_n122_s;
                stage5_col93[3] = fa_s4_c93_n123_s;
                stage5_col93[4] = stage4_col93[6];
                stage5_col94[0] = fa_s4_c93_n122_c;
                stage5_col94[1] = fa_s4_c93_n123_c;
                stage5_col94[2] = fa_s4_c94_n124_s;
                stage5_col94[3] = fa_s4_c94_n125_s;
                stage5_col94[4] = stage4_col94[6];
                stage5_col94[5] = stage4_col94[7];
                stage5_col95[0] = fa_s4_c94_n124_c;
                stage5_col95[1] = fa_s4_c94_n125_c;
                stage5_col95[2] = fa_s4_c95_n126_s;
                stage5_col95[3] = fa_s4_c95_n127_s;
                stage5_col95[4] = stage4_col95[6];
                stage5_col96[0] = fa_s4_c95_n126_c;
                stage5_col96[1] = fa_s4_c95_n127_c;
                stage5_col96[2] = fa_s4_c96_n128_s;
                stage5_col96[3] = fa_s4_c96_n129_s;
                stage5_col96[4] = stage4_col96[6];
                stage5_col96[5] = stage4_col96[7];
                stage5_col97[0] = fa_s4_c96_n128_c;
                stage5_col97[1] = fa_s4_c96_n129_c;
                stage5_col97[2] = fa_s4_c97_n130_s;
                stage5_col97[3] = fa_s4_c97_n131_s;
                stage5_col97[4] = stage4_col97[6];
                stage5_col98[0] = fa_s4_c97_n130_c;
                stage5_col98[1] = fa_s4_c97_n131_c;
                stage5_col98[2] = fa_s4_c98_n132_s;
                stage5_col98[3] = fa_s4_c98_n133_s;
                stage5_col98[4] = stage4_col98[6];
                stage5_col98[5] = stage4_col98[7];
                stage5_col99[0] = fa_s4_c98_n132_c;
                stage5_col99[1] = fa_s4_c98_n133_c;
                stage5_col99[2] = fa_s4_c99_n134_s;
                stage5_col99[3] = fa_s4_c99_n135_s;
                stage5_col99[4] = stage4_col99[6];
                stage5_col100[0] = fa_s4_c99_n134_c;
                stage5_col100[1] = fa_s4_c99_n135_c;
                stage5_col100[2] = fa_s4_c100_n136_s;
                stage5_col100[3] = fa_s4_c100_n137_s;
                stage5_col100[4] = stage4_col100[6];
                stage5_col100[5] = stage4_col100[7];
                stage5_col101[0] = fa_s4_c100_n136_c;
                stage5_col101[1] = fa_s4_c100_n137_c;
                stage5_col101[2] = fa_s4_c101_n138_s;
                stage5_col101[3] = fa_s4_c101_n139_s;
                stage5_col101[4] = stage4_col101[6];
                stage5_col102[0] = fa_s4_c101_n138_c;
                stage5_col102[1] = fa_s4_c101_n139_c;
                stage5_col102[2] = fa_s4_c102_n140_s;
                stage5_col102[3] = fa_s4_c102_n141_s;
                stage5_col102[4] = stage4_col102[6];
                stage5_col102[5] = stage4_col102[7];
                stage5_col103[0] = fa_s4_c102_n140_c;
                stage5_col103[1] = fa_s4_c102_n141_c;
                stage5_col103[2] = fa_s4_c103_n142_s;
                stage5_col103[3] = fa_s4_c103_n143_s;
                stage5_col103[4] = stage4_col103[6];
                stage5_col104[0] = fa_s4_c103_n142_c;
                stage5_col104[1] = fa_s4_c103_n143_c;
                stage5_col104[2] = fa_s4_c104_n144_s;
                stage5_col104[3] = fa_s4_c104_n145_s;
                stage5_col104[4] = stage4_col104[6];
                stage5_col104[5] = stage4_col104[7];
                stage5_col105[0] = fa_s4_c104_n144_c;
                stage5_col105[1] = fa_s4_c104_n145_c;
                stage5_col105[2] = fa_s4_c105_n146_s;
                stage5_col105[3] = fa_s4_c105_n147_s;
                stage5_col105[4] = stage4_col105[6];
                stage5_col106[0] = fa_s4_c105_n146_c;
                stage5_col106[1] = fa_s4_c105_n147_c;
                stage5_col106[2] = fa_s4_c106_n148_s;
                stage5_col106[3] = fa_s4_c106_n149_s;
                stage5_col106[4] = stage4_col106[6];
                stage5_col106[5] = stage4_col106[7];
                stage5_col107[0] = fa_s4_c106_n148_c;
                stage5_col107[1] = fa_s4_c106_n149_c;
                stage5_col107[2] = fa_s4_c107_n150_s;
                stage5_col107[3] = fa_s4_c107_n151_s;
                stage5_col107[4] = stage4_col107[6];
                stage5_col108[0] = fa_s4_c107_n150_c;
                stage5_col108[1] = fa_s4_c107_n151_c;
                stage5_col108[2] = fa_s4_c108_n152_s;
                stage5_col108[3] = fa_s4_c108_n153_s;
                stage5_col108[4] = stage4_col108[6];
                stage5_col108[5] = stage4_col108[7];
                stage5_col109[0] = fa_s4_c108_n152_c;
                stage5_col109[1] = fa_s4_c108_n153_c;
                stage5_col109[2] = fa_s4_c109_n154_s;
                stage5_col109[3] = fa_s4_c109_n155_s;
                stage5_col109[4] = stage4_col109[6];
                stage5_col110[0] = fa_s4_c109_n154_c;
                stage5_col110[1] = fa_s4_c109_n155_c;
                stage5_col110[2] = fa_s4_c110_n156_s;
                stage5_col110[3] = fa_s4_c110_n157_s;
                stage5_col110[4] = stage4_col110[6];
                stage5_col110[5] = stage4_col110[7];
                stage5_col111[0] = fa_s4_c110_n156_c;
                stage5_col111[1] = fa_s4_c110_n157_c;
                stage5_col111[2] = fa_s4_c111_n158_s;
                stage5_col111[3] = fa_s4_c111_n159_s;
                stage5_col111[4] = stage4_col111[6];
                stage5_col112[0] = fa_s4_c111_n158_c;
                stage5_col112[1] = fa_s4_c111_n159_c;
                stage5_col112[2] = fa_s4_c112_n160_s;
                stage5_col112[3] = fa_s4_c112_n161_s;
                stage5_col112[4] = stage4_col112[6];
                stage5_col112[5] = stage4_col112[7];
                stage5_col113[0] = fa_s4_c112_n160_c;
                stage5_col113[1] = fa_s4_c112_n161_c;
                stage5_col113[2] = fa_s4_c113_n162_s;
                stage5_col113[3] = fa_s4_c113_n163_s;
                stage5_col113[4] = stage4_col113[6];
                stage5_col114[0] = fa_s4_c113_n162_c;
                stage5_col114[1] = fa_s4_c113_n163_c;
                stage5_col114[2] = fa_s4_c114_n164_s;
                stage5_col114[3] = fa_s4_c114_n165_s;
                stage5_col114[4] = stage4_col114[6];
                stage5_col114[5] = stage4_col114[7];
                stage5_col115[0] = fa_s4_c114_n164_c;
                stage5_col115[1] = fa_s4_c114_n165_c;
                stage5_col115[2] = fa_s4_c115_n166_s;
                stage5_col115[3] = fa_s4_c115_n167_s;
                stage5_col115[4] = stage4_col115[6];
                stage5_col116[0] = fa_s4_c115_n166_c;
                stage5_col116[1] = fa_s4_c115_n167_c;
                stage5_col116[2] = fa_s4_c116_n168_s;
                stage5_col116[3] = fa_s4_c116_n169_s;
                stage5_col116[4] = stage4_col116[6];
                stage5_col116[5] = stage4_col116[7];
                stage5_col117[0] = fa_s4_c116_n168_c;
                stage5_col117[1] = fa_s4_c116_n169_c;
                stage5_col117[2] = fa_s4_c117_n170_s;
                stage5_col117[3] = fa_s4_c117_n171_s;
                stage5_col117[4] = stage4_col117[6];
                stage5_col118[0] = fa_s4_c117_n170_c;
                stage5_col118[1] = fa_s4_c117_n171_c;
                stage5_col118[2] = fa_s4_c118_n172_s;
                stage5_col118[3] = fa_s4_c118_n173_s;
                stage5_col118[4] = stage4_col118[6];
                stage5_col118[5] = stage4_col118[7];
                stage5_col119[0] = fa_s4_c118_n172_c;
                stage5_col119[1] = fa_s4_c118_n173_c;
                stage5_col119[2] = fa_s4_c119_n174_s;
                stage5_col119[3] = fa_s4_c119_n175_s;
                stage5_col119[4] = stage4_col119[6];
                stage5_col120[0] = fa_s4_c119_n174_c;
                stage5_col120[1] = fa_s4_c119_n175_c;
                stage5_col120[2] = fa_s4_c120_n176_s;
                stage5_col120[3] = fa_s4_c120_n177_s;
                stage5_col120[4] = stage4_col120[6];
                stage5_col120[5] = stage4_col120[7];
                stage5_col121[0] = fa_s4_c120_n176_c;
                stage5_col121[1] = fa_s4_c120_n177_c;
                stage5_col121[2] = fa_s4_c121_n178_s;
                stage5_col121[3] = fa_s4_c121_n179_s;
                stage5_col121[4] = stage4_col121[6];
                stage5_col122[0] = fa_s4_c121_n178_c;
                stage5_col122[1] = fa_s4_c121_n179_c;
                stage5_col122[2] = fa_s4_c122_n180_s;
                stage5_col122[3] = fa_s4_c122_n181_s;
                stage5_col122[4] = stage4_col122[6];
                stage5_col122[5] = stage4_col122[7];
                stage5_col123[0] = fa_s4_c122_n180_c;
                stage5_col123[1] = fa_s4_c122_n181_c;
                stage5_col123[2] = fa_s4_c123_n182_s;
                stage5_col123[3] = fa_s4_c123_n183_s;
                stage5_col123[4] = stage4_col123[6];
                stage5_col124[0] = fa_s4_c123_n182_c;
                stage5_col124[1] = fa_s4_c123_n183_c;
                stage5_col124[2] = fa_s4_c124_n184_s;
                stage5_col124[3] = fa_s4_c124_n185_s;
                stage5_col124[4] = stage4_col124[6];
                stage5_col124[5] = stage4_col124[7];
                stage5_col125[0] = fa_s4_c124_n184_c;
                stage5_col125[1] = fa_s4_c124_n185_c;
                stage5_col125[2] = fa_s4_c125_n186_s;
                stage5_col125[3] = fa_s4_c125_n187_s;
                stage5_col125[4] = stage4_col125[6];
                stage5_col126[0] = fa_s4_c125_n186_c;
                stage5_col126[1] = fa_s4_c125_n187_c;
                stage5_col126[2] = fa_s4_c126_n188_s;
                stage5_col126[3] = fa_s4_c126_n189_s;
                stage5_col126[4] = stage4_col126[6];
                stage5_col126[5] = stage4_col126[7];
                stage5_col127[0] = fa_s4_c126_n188_c;
                stage5_col127[1] = fa_s4_c126_n189_c;
                stage5_col127[2] = stage4_col127[0];
                stage5_col127[3] = stage4_col127[1];
                stage5_col127[4] = stage4_col127[2];
                stage5_col127[5] = stage4_col127[3];
                stage5_col127[6] = stage4_col127[4];
                stage5_col127[7] = stage4_col127[5];
                stage5_col127[8] = stage4_col127[6];
                stage5_col127[9] = stage4_col127[7];
                stage5_col127[10] = stage4_col127[8];
                stage5_col127[11] = stage4_col127[9];
                stage5_col127[12] = stage4_col127[10];
                stage5_col127[13] = stage4_col127[11];
                stage5_col127[14] = stage4_col127[12];
                stage5_col127[15] = stage4_col127[13];
                stage5_col127[16] = stage4_col127[14];
                stage5_col127[17] = stage4_col127[15];
                stage5_col127[18] = stage4_col127[16];
                stage5_col127[19] = stage4_col127[17];
                stage5_col127[20] = stage4_col127[18];
                stage5_col127[21] = stage4_col127[19];
                stage5_col127[22] = stage4_col127[20];
                stage5_col127[23] = stage4_col127[21];
                stage5_col127[24] = stage4_col127[22];
                stage5_col127[25] = stage4_col127[23];
                stage5_col127[26] = stage4_col127[24];
                stage5_col127[27] = stage4_col127[25];
                stage5_col127[28] = stage4_col127[25];
                stage5_col127[29] = stage4_col127[25];
                stage5_col127[30] = stage4_col127[25];
                stage5_col127[31] = stage4_col127[25];
                stage5_col127[32] = stage4_col127[25];
                stage5_col127[33] = stage4_col127[25];
                stage5_col127[34] = stage4_col127[25];
                stage5_col127[35] = stage4_col127[25];
                stage5_col127[36] = stage4_col127[25];
                stage5_col127[37] = stage4_col127[25];
                stage5_col127[38] = stage4_col127[25];
                stage5_col127[39] = stage4_col127[25];
                stage5_col127[40] = stage4_col127[25];
                stage5_col127[41] = stage4_col127[25];
                stage5_col127[42] = stage4_col127[25];
                stage5_col127[43] = stage4_col127[25];
                stage5_col127[44] = stage4_col127[25];
                stage5_col127[45] = stage4_col127[25];
                stage5_col127[46] = stage4_col127[25];
                stage5_col127[47] = stage4_col127[25];
                stage5_col127[48] = stage4_col127[25];
                stage5_col127[49] = stage4_col127[25];
                stage5_col127[50] = stage4_col127[25];
                stage5_col127[51] = stage4_col127[25];
                stage5_col127[52] = stage4_col127[25];
                stage5_col127[53] = stage4_col127[25];
                stage5_col127[54] = stage4_col127[25];
                stage5_col127[55] = stage4_col127[25];
                stage5_col127[56] = stage4_col127[25];
                stage5_col127[57] = stage4_col127[25];
                stage5_col127[58] = stage4_col127[25];
            end
        end
    endgenerate

    // Stage 6: Reduction
    fa fa_s5_c7_n0 (
        .a(stage5_col7[0]),
        .b(stage5_col7[1]),
        .c_in(stage5_col7[2]),
        .s(fa_s5_c7_n0_s),
        .c_out(fa_s5_c7_n0_c)
    );

    fa fa_s5_c28_n1 (
        .a(stage5_col28[0]),
        .b(stage5_col28[1]),
        .c_in(stage5_col28[2]),
        .s(fa_s5_c28_n1_s),
        .c_out(fa_s5_c28_n1_c)
    );

    fa fa_s5_c29_n2 (
        .a(stage5_col29[0]),
        .b(stage5_col29[1]),
        .c_in(stage5_col29[2]),
        .s(fa_s5_c29_n2_s),
        .c_out(fa_s5_c29_n2_c)
    );

    fa fa_s5_c30_n3 (
        .a(stage5_col30[0]),
        .b(stage5_col30[1]),
        .c_in(stage5_col30[2]),
        .s(fa_s5_c30_n3_s),
        .c_out(fa_s5_c30_n3_c)
    );

    fa fa_s5_c31_n4 (
        .a(stage5_col31[0]),
        .b(stage5_col31[1]),
        .c_in(stage5_col31[2]),
        .s(fa_s5_c31_n4_s),
        .c_out(fa_s5_c31_n4_c)
    );

    fa fa_s5_c32_n5 (
        .a(stage5_col32[0]),
        .b(stage5_col32[1]),
        .c_in(stage5_col32[2]),
        .s(fa_s5_c32_n5_s),
        .c_out(fa_s5_c32_n5_c)
    );

    fa fa_s5_c33_n6 (
        .a(stage5_col33[0]),
        .b(stage5_col33[1]),
        .c_in(stage5_col33[2]),
        .s(fa_s5_c33_n6_s),
        .c_out(fa_s5_c33_n6_c)
    );

    fa fa_s5_c34_n7 (
        .a(stage5_col34[0]),
        .b(stage5_col34[1]),
        .c_in(stage5_col34[2]),
        .s(fa_s5_c34_n7_s),
        .c_out(fa_s5_c34_n7_c)
    );

    fa fa_s5_c35_n8 (
        .a(stage5_col35[0]),
        .b(stage5_col35[1]),
        .c_in(stage5_col35[2]),
        .s(fa_s5_c35_n8_s),
        .c_out(fa_s5_c35_n8_c)
    );

    fa fa_s5_c36_n9 (
        .a(stage5_col36[0]),
        .b(stage5_col36[1]),
        .c_in(stage5_col36[2]),
        .s(fa_s5_c36_n9_s),
        .c_out(fa_s5_c36_n9_c)
    );

    fa fa_s5_c37_n10 (
        .a(stage5_col37[0]),
        .b(stage5_col37[1]),
        .c_in(stage5_col37[2]),
        .s(fa_s5_c37_n10_s),
        .c_out(fa_s5_c37_n10_c)
    );

    fa fa_s5_c38_n11 (
        .a(stage5_col38[0]),
        .b(stage5_col38[1]),
        .c_in(stage5_col38[2]),
        .s(fa_s5_c38_n11_s),
        .c_out(fa_s5_c38_n11_c)
    );

    fa fa_s5_c39_n12 (
        .a(stage5_col39[0]),
        .b(stage5_col39[1]),
        .c_in(stage5_col39[2]),
        .s(fa_s5_c39_n12_s),
        .c_out(fa_s5_c39_n12_c)
    );

    fa fa_s5_c40_n13 (
        .a(stage5_col40[0]),
        .b(stage5_col40[1]),
        .c_in(stage5_col40[2]),
        .s(fa_s5_c40_n13_s),
        .c_out(fa_s5_c40_n13_c)
    );

    fa fa_s5_c41_n14 (
        .a(stage5_col41[0]),
        .b(stage5_col41[1]),
        .c_in(stage5_col41[2]),
        .s(fa_s5_c41_n14_s),
        .c_out(fa_s5_c41_n14_c)
    );

    fa fa_s5_c42_n15 (
        .a(stage5_col42[0]),
        .b(stage5_col42[1]),
        .c_in(stage5_col42[2]),
        .s(fa_s5_c42_n15_s),
        .c_out(fa_s5_c42_n15_c)
    );

    fa fa_s5_c43_n16 (
        .a(stage5_col43[0]),
        .b(stage5_col43[1]),
        .c_in(stage5_col43[2]),
        .s(fa_s5_c43_n16_s),
        .c_out(fa_s5_c43_n16_c)
    );

    fa fa_s5_c44_n17 (
        .a(stage5_col44[0]),
        .b(stage5_col44[1]),
        .c_in(stage5_col44[2]),
        .s(fa_s5_c44_n17_s),
        .c_out(fa_s5_c44_n17_c)
    );

    fa fa_s5_c45_n18 (
        .a(stage5_col45[0]),
        .b(stage5_col45[1]),
        .c_in(stage5_col45[2]),
        .s(fa_s5_c45_n18_s),
        .c_out(fa_s5_c45_n18_c)
    );

    fa fa_s5_c46_n19 (
        .a(stage5_col46[0]),
        .b(stage5_col46[1]),
        .c_in(stage5_col46[2]),
        .s(fa_s5_c46_n19_s),
        .c_out(fa_s5_c46_n19_c)
    );

    fa fa_s5_c47_n20 (
        .a(stage5_col47[0]),
        .b(stage5_col47[1]),
        .c_in(stage5_col47[2]),
        .s(fa_s5_c47_n20_s),
        .c_out(fa_s5_c47_n20_c)
    );

    fa fa_s5_c48_n21 (
        .a(stage5_col48[0]),
        .b(stage5_col48[1]),
        .c_in(stage5_col48[2]),
        .s(fa_s5_c48_n21_s),
        .c_out(fa_s5_c48_n21_c)
    );

    fa fa_s5_c49_n22 (
        .a(stage5_col49[0]),
        .b(stage5_col49[1]),
        .c_in(stage5_col49[2]),
        .s(fa_s5_c49_n22_s),
        .c_out(fa_s5_c49_n22_c)
    );

    fa fa_s5_c50_n23 (
        .a(stage5_col50[0]),
        .b(stage5_col50[1]),
        .c_in(stage5_col50[2]),
        .s(fa_s5_c50_n23_s),
        .c_out(fa_s5_c50_n23_c)
    );

    fa fa_s5_c51_n24 (
        .a(stage5_col51[0]),
        .b(stage5_col51[1]),
        .c_in(stage5_col51[2]),
        .s(fa_s5_c51_n24_s),
        .c_out(fa_s5_c51_n24_c)
    );

    fa fa_s5_c52_n25 (
        .a(stage5_col52[0]),
        .b(stage5_col52[1]),
        .c_in(stage5_col52[2]),
        .s(fa_s5_c52_n25_s),
        .c_out(fa_s5_c52_n25_c)
    );

    fa fa_s5_c53_n26 (
        .a(stage5_col53[0]),
        .b(stage5_col53[1]),
        .c_in(stage5_col53[2]),
        .s(fa_s5_c53_n26_s),
        .c_out(fa_s5_c53_n26_c)
    );

    fa fa_s5_c54_n27 (
        .a(stage5_col54[0]),
        .b(stage5_col54[1]),
        .c_in(stage5_col54[2]),
        .s(fa_s5_c54_n27_s),
        .c_out(fa_s5_c54_n27_c)
    );

    fa fa_s5_c55_n28 (
        .a(stage5_col55[0]),
        .b(stage5_col55[1]),
        .c_in(stage5_col55[2]),
        .s(fa_s5_c55_n28_s),
        .c_out(fa_s5_c55_n28_c)
    );

    fa fa_s5_c56_n29 (
        .a(stage5_col56[0]),
        .b(stage5_col56[1]),
        .c_in(stage5_col56[2]),
        .s(fa_s5_c56_n29_s),
        .c_out(fa_s5_c56_n29_c)
    );

    fa fa_s5_c57_n30 (
        .a(stage5_col57[0]),
        .b(stage5_col57[1]),
        .c_in(stage5_col57[2]),
        .s(fa_s5_c57_n30_s),
        .c_out(fa_s5_c57_n30_c)
    );

    fa fa_s5_c58_n31 (
        .a(stage5_col58[0]),
        .b(stage5_col58[1]),
        .c_in(stage5_col58[2]),
        .s(fa_s5_c58_n31_s),
        .c_out(fa_s5_c58_n31_c)
    );

    fa fa_s5_c59_n32 (
        .a(stage5_col59[0]),
        .b(stage5_col59[1]),
        .c_in(stage5_col59[2]),
        .s(fa_s5_c59_n32_s),
        .c_out(fa_s5_c59_n32_c)
    );

    fa fa_s5_c59_n33 (
        .a(stage5_col59[3]),
        .b(stage5_col59[4]),
        .c_in(stage5_col59[5]),
        .s(fa_s5_c59_n33_s),
        .c_out(fa_s5_c59_n33_c)
    );

    fa fa_s5_c60_n34 (
        .a(stage5_col60[0]),
        .b(stage5_col60[1]),
        .c_in(stage5_col60[2]),
        .s(fa_s5_c60_n34_s),
        .c_out(fa_s5_c60_n34_c)
    );

    fa fa_s5_c61_n35 (
        .a(stage5_col61[0]),
        .b(stage5_col61[1]),
        .c_in(stage5_col61[2]),
        .s(fa_s5_c61_n35_s),
        .c_out(fa_s5_c61_n35_c)
    );

    fa fa_s5_c62_n36 (
        .a(stage5_col62[0]),
        .b(stage5_col62[1]),
        .c_in(stage5_col62[2]),
        .s(fa_s5_c62_n36_s),
        .c_out(fa_s5_c62_n36_c)
    );

    fa fa_s5_c63_n37 (
        .a(stage5_col63[0]),
        .b(stage5_col63[1]),
        .c_in(stage5_col63[2]),
        .s(fa_s5_c63_n37_s),
        .c_out(fa_s5_c63_n37_c)
    );

    fa fa_s5_c64_n38 (
        .a(stage5_col64[0]),
        .b(stage5_col64[1]),
        .c_in(stage5_col64[2]),
        .s(fa_s5_c64_n38_s),
        .c_out(fa_s5_c64_n38_c)
    );

    fa fa_s5_c64_n39 (
        .a(stage5_col64[3]),
        .b(stage5_col64[4]),
        .c_in(stage5_col64[5]),
        .s(fa_s5_c64_n39_s),
        .c_out(fa_s5_c64_n39_c)
    );

    fa fa_s5_c65_n40 (
        .a(stage5_col65[0]),
        .b(stage5_col65[1]),
        .c_in(stage5_col65[2]),
        .s(fa_s5_c65_n40_s),
        .c_out(fa_s5_c65_n40_c)
    );

    fa fa_s5_c66_n41 (
        .a(stage5_col66[0]),
        .b(stage5_col66[1]),
        .c_in(stage5_col66[2]),
        .s(fa_s5_c66_n41_s),
        .c_out(fa_s5_c66_n41_c)
    );

    fa fa_s5_c66_n42 (
        .a(stage5_col66[3]),
        .b(stage5_col66[4]),
        .c_in(stage5_col66[5]),
        .s(fa_s5_c66_n42_s),
        .c_out(fa_s5_c66_n42_c)
    );

    fa fa_s5_c67_n43 (
        .a(stage5_col67[0]),
        .b(stage5_col67[1]),
        .c_in(stage5_col67[2]),
        .s(fa_s5_c67_n43_s),
        .c_out(fa_s5_c67_n43_c)
    );

    fa fa_s5_c68_n44 (
        .a(stage5_col68[0]),
        .b(stage5_col68[1]),
        .c_in(stage5_col68[2]),
        .s(fa_s5_c68_n44_s),
        .c_out(fa_s5_c68_n44_c)
    );

    fa fa_s5_c68_n45 (
        .a(stage5_col68[3]),
        .b(stage5_col68[4]),
        .c_in(stage5_col68[5]),
        .s(fa_s5_c68_n45_s),
        .c_out(fa_s5_c68_n45_c)
    );

    fa fa_s5_c69_n46 (
        .a(stage5_col69[0]),
        .b(stage5_col69[1]),
        .c_in(stage5_col69[2]),
        .s(fa_s5_c69_n46_s),
        .c_out(fa_s5_c69_n46_c)
    );

    fa fa_s5_c70_n47 (
        .a(stage5_col70[0]),
        .b(stage5_col70[1]),
        .c_in(stage5_col70[2]),
        .s(fa_s5_c70_n47_s),
        .c_out(fa_s5_c70_n47_c)
    );

    fa fa_s5_c70_n48 (
        .a(stage5_col70[3]),
        .b(stage5_col70[4]),
        .c_in(stage5_col70[5]),
        .s(fa_s5_c70_n48_s),
        .c_out(fa_s5_c70_n48_c)
    );

    fa fa_s5_c71_n49 (
        .a(stage5_col71[0]),
        .b(stage5_col71[1]),
        .c_in(stage5_col71[2]),
        .s(fa_s5_c71_n49_s),
        .c_out(fa_s5_c71_n49_c)
    );

    fa fa_s5_c72_n50 (
        .a(stage5_col72[0]),
        .b(stage5_col72[1]),
        .c_in(stage5_col72[2]),
        .s(fa_s5_c72_n50_s),
        .c_out(fa_s5_c72_n50_c)
    );

    fa fa_s5_c72_n51 (
        .a(stage5_col72[3]),
        .b(stage5_col72[4]),
        .c_in(stage5_col72[5]),
        .s(fa_s5_c72_n51_s),
        .c_out(fa_s5_c72_n51_c)
    );

    fa fa_s5_c73_n52 (
        .a(stage5_col73[0]),
        .b(stage5_col73[1]),
        .c_in(stage5_col73[2]),
        .s(fa_s5_c73_n52_s),
        .c_out(fa_s5_c73_n52_c)
    );

    fa fa_s5_c74_n53 (
        .a(stage5_col74[0]),
        .b(stage5_col74[1]),
        .c_in(stage5_col74[2]),
        .s(fa_s5_c74_n53_s),
        .c_out(fa_s5_c74_n53_c)
    );

    fa fa_s5_c74_n54 (
        .a(stage5_col74[3]),
        .b(stage5_col74[4]),
        .c_in(stage5_col74[5]),
        .s(fa_s5_c74_n54_s),
        .c_out(fa_s5_c74_n54_c)
    );

    fa fa_s5_c75_n55 (
        .a(stage5_col75[0]),
        .b(stage5_col75[1]),
        .c_in(stage5_col75[2]),
        .s(fa_s5_c75_n55_s),
        .c_out(fa_s5_c75_n55_c)
    );

    fa fa_s5_c76_n56 (
        .a(stage5_col76[0]),
        .b(stage5_col76[1]),
        .c_in(stage5_col76[2]),
        .s(fa_s5_c76_n56_s),
        .c_out(fa_s5_c76_n56_c)
    );

    fa fa_s5_c76_n57 (
        .a(stage5_col76[3]),
        .b(stage5_col76[4]),
        .c_in(stage5_col76[5]),
        .s(fa_s5_c76_n57_s),
        .c_out(fa_s5_c76_n57_c)
    );

    fa fa_s5_c77_n58 (
        .a(stage5_col77[0]),
        .b(stage5_col77[1]),
        .c_in(stage5_col77[2]),
        .s(fa_s5_c77_n58_s),
        .c_out(fa_s5_c77_n58_c)
    );

    fa fa_s5_c78_n59 (
        .a(stage5_col78[0]),
        .b(stage5_col78[1]),
        .c_in(stage5_col78[2]),
        .s(fa_s5_c78_n59_s),
        .c_out(fa_s5_c78_n59_c)
    );

    fa fa_s5_c78_n60 (
        .a(stage5_col78[3]),
        .b(stage5_col78[4]),
        .c_in(stage5_col78[5]),
        .s(fa_s5_c78_n60_s),
        .c_out(fa_s5_c78_n60_c)
    );

    fa fa_s5_c79_n61 (
        .a(stage5_col79[0]),
        .b(stage5_col79[1]),
        .c_in(stage5_col79[2]),
        .s(fa_s5_c79_n61_s),
        .c_out(fa_s5_c79_n61_c)
    );

    fa fa_s5_c80_n62 (
        .a(stage5_col80[0]),
        .b(stage5_col80[1]),
        .c_in(stage5_col80[2]),
        .s(fa_s5_c80_n62_s),
        .c_out(fa_s5_c80_n62_c)
    );

    fa fa_s5_c80_n63 (
        .a(stage5_col80[3]),
        .b(stage5_col80[4]),
        .c_in(stage5_col80[5]),
        .s(fa_s5_c80_n63_s),
        .c_out(fa_s5_c80_n63_c)
    );

    fa fa_s5_c81_n64 (
        .a(stage5_col81[0]),
        .b(stage5_col81[1]),
        .c_in(stage5_col81[2]),
        .s(fa_s5_c81_n64_s),
        .c_out(fa_s5_c81_n64_c)
    );

    fa fa_s5_c82_n65 (
        .a(stage5_col82[0]),
        .b(stage5_col82[1]),
        .c_in(stage5_col82[2]),
        .s(fa_s5_c82_n65_s),
        .c_out(fa_s5_c82_n65_c)
    );

    fa fa_s5_c82_n66 (
        .a(stage5_col82[3]),
        .b(stage5_col82[4]),
        .c_in(stage5_col82[5]),
        .s(fa_s5_c82_n66_s),
        .c_out(fa_s5_c82_n66_c)
    );

    fa fa_s5_c83_n67 (
        .a(stage5_col83[0]),
        .b(stage5_col83[1]),
        .c_in(stage5_col83[2]),
        .s(fa_s5_c83_n67_s),
        .c_out(fa_s5_c83_n67_c)
    );

    fa fa_s5_c84_n68 (
        .a(stage5_col84[0]),
        .b(stage5_col84[1]),
        .c_in(stage5_col84[2]),
        .s(fa_s5_c84_n68_s),
        .c_out(fa_s5_c84_n68_c)
    );

    fa fa_s5_c84_n69 (
        .a(stage5_col84[3]),
        .b(stage5_col84[4]),
        .c_in(stage5_col84[5]),
        .s(fa_s5_c84_n69_s),
        .c_out(fa_s5_c84_n69_c)
    );

    fa fa_s5_c85_n70 (
        .a(stage5_col85[0]),
        .b(stage5_col85[1]),
        .c_in(stage5_col85[2]),
        .s(fa_s5_c85_n70_s),
        .c_out(fa_s5_c85_n70_c)
    );

    fa fa_s5_c86_n71 (
        .a(stage5_col86[0]),
        .b(stage5_col86[1]),
        .c_in(stage5_col86[2]),
        .s(fa_s5_c86_n71_s),
        .c_out(fa_s5_c86_n71_c)
    );

    fa fa_s5_c86_n72 (
        .a(stage5_col86[3]),
        .b(stage5_col86[4]),
        .c_in(stage5_col86[5]),
        .s(fa_s5_c86_n72_s),
        .c_out(fa_s5_c86_n72_c)
    );

    fa fa_s5_c87_n73 (
        .a(stage5_col87[0]),
        .b(stage5_col87[1]),
        .c_in(stage5_col87[2]),
        .s(fa_s5_c87_n73_s),
        .c_out(fa_s5_c87_n73_c)
    );

    fa fa_s5_c88_n74 (
        .a(stage5_col88[0]),
        .b(stage5_col88[1]),
        .c_in(stage5_col88[2]),
        .s(fa_s5_c88_n74_s),
        .c_out(fa_s5_c88_n74_c)
    );

    fa fa_s5_c88_n75 (
        .a(stage5_col88[3]),
        .b(stage5_col88[4]),
        .c_in(stage5_col88[5]),
        .s(fa_s5_c88_n75_s),
        .c_out(fa_s5_c88_n75_c)
    );

    fa fa_s5_c89_n76 (
        .a(stage5_col89[0]),
        .b(stage5_col89[1]),
        .c_in(stage5_col89[2]),
        .s(fa_s5_c89_n76_s),
        .c_out(fa_s5_c89_n76_c)
    );

    fa fa_s5_c90_n77 (
        .a(stage5_col90[0]),
        .b(stage5_col90[1]),
        .c_in(stage5_col90[2]),
        .s(fa_s5_c90_n77_s),
        .c_out(fa_s5_c90_n77_c)
    );

    fa fa_s5_c90_n78 (
        .a(stage5_col90[3]),
        .b(stage5_col90[4]),
        .c_in(stage5_col90[5]),
        .s(fa_s5_c90_n78_s),
        .c_out(fa_s5_c90_n78_c)
    );

    fa fa_s5_c91_n79 (
        .a(stage5_col91[0]),
        .b(stage5_col91[1]),
        .c_in(stage5_col91[2]),
        .s(fa_s5_c91_n79_s),
        .c_out(fa_s5_c91_n79_c)
    );

    fa fa_s5_c92_n80 (
        .a(stage5_col92[0]),
        .b(stage5_col92[1]),
        .c_in(stage5_col92[2]),
        .s(fa_s5_c92_n80_s),
        .c_out(fa_s5_c92_n80_c)
    );

    fa fa_s5_c92_n81 (
        .a(stage5_col92[3]),
        .b(stage5_col92[4]),
        .c_in(stage5_col92[5]),
        .s(fa_s5_c92_n81_s),
        .c_out(fa_s5_c92_n81_c)
    );

    fa fa_s5_c93_n82 (
        .a(stage5_col93[0]),
        .b(stage5_col93[1]),
        .c_in(stage5_col93[2]),
        .s(fa_s5_c93_n82_s),
        .c_out(fa_s5_c93_n82_c)
    );

    fa fa_s5_c94_n83 (
        .a(stage5_col94[0]),
        .b(stage5_col94[1]),
        .c_in(stage5_col94[2]),
        .s(fa_s5_c94_n83_s),
        .c_out(fa_s5_c94_n83_c)
    );

    fa fa_s5_c94_n84 (
        .a(stage5_col94[3]),
        .b(stage5_col94[4]),
        .c_in(stage5_col94[5]),
        .s(fa_s5_c94_n84_s),
        .c_out(fa_s5_c94_n84_c)
    );

    fa fa_s5_c95_n85 (
        .a(stage5_col95[0]),
        .b(stage5_col95[1]),
        .c_in(stage5_col95[2]),
        .s(fa_s5_c95_n85_s),
        .c_out(fa_s5_c95_n85_c)
    );

    fa fa_s5_c96_n86 (
        .a(stage5_col96[0]),
        .b(stage5_col96[1]),
        .c_in(stage5_col96[2]),
        .s(fa_s5_c96_n86_s),
        .c_out(fa_s5_c96_n86_c)
    );

    fa fa_s5_c96_n87 (
        .a(stage5_col96[3]),
        .b(stage5_col96[4]),
        .c_in(stage5_col96[5]),
        .s(fa_s5_c96_n87_s),
        .c_out(fa_s5_c96_n87_c)
    );

    fa fa_s5_c97_n88 (
        .a(stage5_col97[0]),
        .b(stage5_col97[1]),
        .c_in(stage5_col97[2]),
        .s(fa_s5_c97_n88_s),
        .c_out(fa_s5_c97_n88_c)
    );

    fa fa_s5_c98_n89 (
        .a(stage5_col98[0]),
        .b(stage5_col98[1]),
        .c_in(stage5_col98[2]),
        .s(fa_s5_c98_n89_s),
        .c_out(fa_s5_c98_n89_c)
    );

    fa fa_s5_c98_n90 (
        .a(stage5_col98[3]),
        .b(stage5_col98[4]),
        .c_in(stage5_col98[5]),
        .s(fa_s5_c98_n90_s),
        .c_out(fa_s5_c98_n90_c)
    );

    fa fa_s5_c99_n91 (
        .a(stage5_col99[0]),
        .b(stage5_col99[1]),
        .c_in(stage5_col99[2]),
        .s(fa_s5_c99_n91_s),
        .c_out(fa_s5_c99_n91_c)
    );

    fa fa_s5_c100_n92 (
        .a(stage5_col100[0]),
        .b(stage5_col100[1]),
        .c_in(stage5_col100[2]),
        .s(fa_s5_c100_n92_s),
        .c_out(fa_s5_c100_n92_c)
    );

    fa fa_s5_c100_n93 (
        .a(stage5_col100[3]),
        .b(stage5_col100[4]),
        .c_in(stage5_col100[5]),
        .s(fa_s5_c100_n93_s),
        .c_out(fa_s5_c100_n93_c)
    );

    fa fa_s5_c101_n94 (
        .a(stage5_col101[0]),
        .b(stage5_col101[1]),
        .c_in(stage5_col101[2]),
        .s(fa_s5_c101_n94_s),
        .c_out(fa_s5_c101_n94_c)
    );

    fa fa_s5_c102_n95 (
        .a(stage5_col102[0]),
        .b(stage5_col102[1]),
        .c_in(stage5_col102[2]),
        .s(fa_s5_c102_n95_s),
        .c_out(fa_s5_c102_n95_c)
    );

    fa fa_s5_c102_n96 (
        .a(stage5_col102[3]),
        .b(stage5_col102[4]),
        .c_in(stage5_col102[5]),
        .s(fa_s5_c102_n96_s),
        .c_out(fa_s5_c102_n96_c)
    );

    fa fa_s5_c103_n97 (
        .a(stage5_col103[0]),
        .b(stage5_col103[1]),
        .c_in(stage5_col103[2]),
        .s(fa_s5_c103_n97_s),
        .c_out(fa_s5_c103_n97_c)
    );

    fa fa_s5_c104_n98 (
        .a(stage5_col104[0]),
        .b(stage5_col104[1]),
        .c_in(stage5_col104[2]),
        .s(fa_s5_c104_n98_s),
        .c_out(fa_s5_c104_n98_c)
    );

    fa fa_s5_c104_n99 (
        .a(stage5_col104[3]),
        .b(stage5_col104[4]),
        .c_in(stage5_col104[5]),
        .s(fa_s5_c104_n99_s),
        .c_out(fa_s5_c104_n99_c)
    );

    fa fa_s5_c105_n100 (
        .a(stage5_col105[0]),
        .b(stage5_col105[1]),
        .c_in(stage5_col105[2]),
        .s(fa_s5_c105_n100_s),
        .c_out(fa_s5_c105_n100_c)
    );

    fa fa_s5_c106_n101 (
        .a(stage5_col106[0]),
        .b(stage5_col106[1]),
        .c_in(stage5_col106[2]),
        .s(fa_s5_c106_n101_s),
        .c_out(fa_s5_c106_n101_c)
    );

    fa fa_s5_c106_n102 (
        .a(stage5_col106[3]),
        .b(stage5_col106[4]),
        .c_in(stage5_col106[5]),
        .s(fa_s5_c106_n102_s),
        .c_out(fa_s5_c106_n102_c)
    );

    fa fa_s5_c107_n103 (
        .a(stage5_col107[0]),
        .b(stage5_col107[1]),
        .c_in(stage5_col107[2]),
        .s(fa_s5_c107_n103_s),
        .c_out(fa_s5_c107_n103_c)
    );

    fa fa_s5_c108_n104 (
        .a(stage5_col108[0]),
        .b(stage5_col108[1]),
        .c_in(stage5_col108[2]),
        .s(fa_s5_c108_n104_s),
        .c_out(fa_s5_c108_n104_c)
    );

    fa fa_s5_c108_n105 (
        .a(stage5_col108[3]),
        .b(stage5_col108[4]),
        .c_in(stage5_col108[5]),
        .s(fa_s5_c108_n105_s),
        .c_out(fa_s5_c108_n105_c)
    );

    fa fa_s5_c109_n106 (
        .a(stage5_col109[0]),
        .b(stage5_col109[1]),
        .c_in(stage5_col109[2]),
        .s(fa_s5_c109_n106_s),
        .c_out(fa_s5_c109_n106_c)
    );

    fa fa_s5_c110_n107 (
        .a(stage5_col110[0]),
        .b(stage5_col110[1]),
        .c_in(stage5_col110[2]),
        .s(fa_s5_c110_n107_s),
        .c_out(fa_s5_c110_n107_c)
    );

    fa fa_s5_c110_n108 (
        .a(stage5_col110[3]),
        .b(stage5_col110[4]),
        .c_in(stage5_col110[5]),
        .s(fa_s5_c110_n108_s),
        .c_out(fa_s5_c110_n108_c)
    );

    fa fa_s5_c111_n109 (
        .a(stage5_col111[0]),
        .b(stage5_col111[1]),
        .c_in(stage5_col111[2]),
        .s(fa_s5_c111_n109_s),
        .c_out(fa_s5_c111_n109_c)
    );

    fa fa_s5_c112_n110 (
        .a(stage5_col112[0]),
        .b(stage5_col112[1]),
        .c_in(stage5_col112[2]),
        .s(fa_s5_c112_n110_s),
        .c_out(fa_s5_c112_n110_c)
    );

    fa fa_s5_c112_n111 (
        .a(stage5_col112[3]),
        .b(stage5_col112[4]),
        .c_in(stage5_col112[5]),
        .s(fa_s5_c112_n111_s),
        .c_out(fa_s5_c112_n111_c)
    );

    fa fa_s5_c113_n112 (
        .a(stage5_col113[0]),
        .b(stage5_col113[1]),
        .c_in(stage5_col113[2]),
        .s(fa_s5_c113_n112_s),
        .c_out(fa_s5_c113_n112_c)
    );

    fa fa_s5_c114_n113 (
        .a(stage5_col114[0]),
        .b(stage5_col114[1]),
        .c_in(stage5_col114[2]),
        .s(fa_s5_c114_n113_s),
        .c_out(fa_s5_c114_n113_c)
    );

    fa fa_s5_c114_n114 (
        .a(stage5_col114[3]),
        .b(stage5_col114[4]),
        .c_in(stage5_col114[5]),
        .s(fa_s5_c114_n114_s),
        .c_out(fa_s5_c114_n114_c)
    );

    fa fa_s5_c115_n115 (
        .a(stage5_col115[0]),
        .b(stage5_col115[1]),
        .c_in(stage5_col115[2]),
        .s(fa_s5_c115_n115_s),
        .c_out(fa_s5_c115_n115_c)
    );

    fa fa_s5_c116_n116 (
        .a(stage5_col116[0]),
        .b(stage5_col116[1]),
        .c_in(stage5_col116[2]),
        .s(fa_s5_c116_n116_s),
        .c_out(fa_s5_c116_n116_c)
    );

    fa fa_s5_c116_n117 (
        .a(stage5_col116[3]),
        .b(stage5_col116[4]),
        .c_in(stage5_col116[5]),
        .s(fa_s5_c116_n117_s),
        .c_out(fa_s5_c116_n117_c)
    );

    fa fa_s5_c117_n118 (
        .a(stage5_col117[0]),
        .b(stage5_col117[1]),
        .c_in(stage5_col117[2]),
        .s(fa_s5_c117_n118_s),
        .c_out(fa_s5_c117_n118_c)
    );

    fa fa_s5_c118_n119 (
        .a(stage5_col118[0]),
        .b(stage5_col118[1]),
        .c_in(stage5_col118[2]),
        .s(fa_s5_c118_n119_s),
        .c_out(fa_s5_c118_n119_c)
    );

    fa fa_s5_c118_n120 (
        .a(stage5_col118[3]),
        .b(stage5_col118[4]),
        .c_in(stage5_col118[5]),
        .s(fa_s5_c118_n120_s),
        .c_out(fa_s5_c118_n120_c)
    );

    fa fa_s5_c119_n121 (
        .a(stage5_col119[0]),
        .b(stage5_col119[1]),
        .c_in(stage5_col119[2]),
        .s(fa_s5_c119_n121_s),
        .c_out(fa_s5_c119_n121_c)
    );

    fa fa_s5_c120_n122 (
        .a(stage5_col120[0]),
        .b(stage5_col120[1]),
        .c_in(stage5_col120[2]),
        .s(fa_s5_c120_n122_s),
        .c_out(fa_s5_c120_n122_c)
    );

    fa fa_s5_c120_n123 (
        .a(stage5_col120[3]),
        .b(stage5_col120[4]),
        .c_in(stage5_col120[5]),
        .s(fa_s5_c120_n123_s),
        .c_out(fa_s5_c120_n123_c)
    );

    fa fa_s5_c121_n124 (
        .a(stage5_col121[0]),
        .b(stage5_col121[1]),
        .c_in(stage5_col121[2]),
        .s(fa_s5_c121_n124_s),
        .c_out(fa_s5_c121_n124_c)
    );

    fa fa_s5_c122_n125 (
        .a(stage5_col122[0]),
        .b(stage5_col122[1]),
        .c_in(stage5_col122[2]),
        .s(fa_s5_c122_n125_s),
        .c_out(fa_s5_c122_n125_c)
    );

    fa fa_s5_c122_n126 (
        .a(stage5_col122[3]),
        .b(stage5_col122[4]),
        .c_in(stage5_col122[5]),
        .s(fa_s5_c122_n126_s),
        .c_out(fa_s5_c122_n126_c)
    );

    fa fa_s5_c123_n127 (
        .a(stage5_col123[0]),
        .b(stage5_col123[1]),
        .c_in(stage5_col123[2]),
        .s(fa_s5_c123_n127_s),
        .c_out(fa_s5_c123_n127_c)
    );

    fa fa_s5_c124_n128 (
        .a(stage5_col124[0]),
        .b(stage5_col124[1]),
        .c_in(stage5_col124[2]),
        .s(fa_s5_c124_n128_s),
        .c_out(fa_s5_c124_n128_c)
    );

    fa fa_s5_c124_n129 (
        .a(stage5_col124[3]),
        .b(stage5_col124[4]),
        .c_in(stage5_col124[5]),
        .s(fa_s5_c124_n129_s),
        .c_out(fa_s5_c124_n129_c)
    );

    fa fa_s5_c125_n130 (
        .a(stage5_col125[0]),
        .b(stage5_col125[1]),
        .c_in(stage5_col125[2]),
        .s(fa_s5_c125_n130_s),
        .c_out(fa_s5_c125_n130_c)
    );

    fa fa_s5_c126_n131 (
        .a(stage5_col126[0]),
        .b(stage5_col126[1]),
        .c_in(stage5_col126[2]),
        .s(fa_s5_c126_n131_s),
        .c_out(fa_s5_c126_n131_c)
    );

    fa fa_s5_c126_n132 (
        .a(stage5_col126[3]),
        .b(stage5_col126[4]),
        .c_in(stage5_col126[5]),
        .s(fa_s5_c126_n132_s),
        .c_out(fa_s5_c126_n132_c)
    );

    ha ha_s5_c5_n0 (
        .a(stage5_col5[0]),
        .b(stage5_col5[1]),
        .s(ha_s5_c5_n0_s),
        .c_out(ha_s5_c5_n0_c)
    );

    ha ha_s5_c60_n1 (
        .a(stage5_col60[3]),
        .b(stage5_col60[4]),
        .s(ha_s5_c60_n1_s),
        .c_out(ha_s5_c60_n1_c)
    );

    ha ha_s5_c61_n2 (
        .a(stage5_col61[3]),
        .b(stage5_col61[4]),
        .s(ha_s5_c61_n2_s),
        .c_out(ha_s5_c61_n2_c)
    );

    ha ha_s5_c62_n3 (
        .a(stage5_col62[3]),
        .b(stage5_col62[4]),
        .s(ha_s5_c62_n3_s),
        .c_out(ha_s5_c62_n3_c)
    );

    ha ha_s5_c63_n4 (
        .a(stage5_col63[3]),
        .b(stage5_col63[4]),
        .s(ha_s5_c63_n4_s),
        .c_out(ha_s5_c63_n4_c)
    );

    ha ha_s5_c65_n5 (
        .a(stage5_col65[3]),
        .b(stage5_col65[4]),
        .s(ha_s5_c65_n5_s),
        .c_out(ha_s5_c65_n5_c)
    );

    ha ha_s5_c67_n6 (
        .a(stage5_col67[3]),
        .b(stage5_col67[4]),
        .s(ha_s5_c67_n6_s),
        .c_out(ha_s5_c67_n6_c)
    );

    ha ha_s5_c69_n7 (
        .a(stage5_col69[3]),
        .b(stage5_col69[4]),
        .s(ha_s5_c69_n7_s),
        .c_out(ha_s5_c69_n7_c)
    );

    ha ha_s5_c71_n8 (
        .a(stage5_col71[3]),
        .b(stage5_col71[4]),
        .s(ha_s5_c71_n8_s),
        .c_out(ha_s5_c71_n8_c)
    );

    ha ha_s5_c73_n9 (
        .a(stage5_col73[3]),
        .b(stage5_col73[4]),
        .s(ha_s5_c73_n9_s),
        .c_out(ha_s5_c73_n9_c)
    );

    ha ha_s5_c75_n10 (
        .a(stage5_col75[3]),
        .b(stage5_col75[4]),
        .s(ha_s5_c75_n10_s),
        .c_out(ha_s5_c75_n10_c)
    );

    ha ha_s5_c77_n11 (
        .a(stage5_col77[3]),
        .b(stage5_col77[4]),
        .s(ha_s5_c77_n11_s),
        .c_out(ha_s5_c77_n11_c)
    );

    ha ha_s5_c79_n12 (
        .a(stage5_col79[3]),
        .b(stage5_col79[4]),
        .s(ha_s5_c79_n12_s),
        .c_out(ha_s5_c79_n12_c)
    );

    ha ha_s5_c81_n13 (
        .a(stage5_col81[3]),
        .b(stage5_col81[4]),
        .s(ha_s5_c81_n13_s),
        .c_out(ha_s5_c81_n13_c)
    );

    ha ha_s5_c83_n14 (
        .a(stage5_col83[3]),
        .b(stage5_col83[4]),
        .s(ha_s5_c83_n14_s),
        .c_out(ha_s5_c83_n14_c)
    );

    ha ha_s5_c85_n15 (
        .a(stage5_col85[3]),
        .b(stage5_col85[4]),
        .s(ha_s5_c85_n15_s),
        .c_out(ha_s5_c85_n15_c)
    );

    ha ha_s5_c87_n16 (
        .a(stage5_col87[3]),
        .b(stage5_col87[4]),
        .s(ha_s5_c87_n16_s),
        .c_out(ha_s5_c87_n16_c)
    );

    ha ha_s5_c89_n17 (
        .a(stage5_col89[3]),
        .b(stage5_col89[4]),
        .s(ha_s5_c89_n17_s),
        .c_out(ha_s5_c89_n17_c)
    );

    ha ha_s5_c91_n18 (
        .a(stage5_col91[3]),
        .b(stage5_col91[4]),
        .s(ha_s5_c91_n18_s),
        .c_out(ha_s5_c91_n18_c)
    );

    ha ha_s5_c93_n19 (
        .a(stage5_col93[3]),
        .b(stage5_col93[4]),
        .s(ha_s5_c93_n19_s),
        .c_out(ha_s5_c93_n19_c)
    );

    ha ha_s5_c95_n20 (
        .a(stage5_col95[3]),
        .b(stage5_col95[4]),
        .s(ha_s5_c95_n20_s),
        .c_out(ha_s5_c95_n20_c)
    );

    ha ha_s5_c97_n21 (
        .a(stage5_col97[3]),
        .b(stage5_col97[4]),
        .s(ha_s5_c97_n21_s),
        .c_out(ha_s5_c97_n21_c)
    );

    ha ha_s5_c99_n22 (
        .a(stage5_col99[3]),
        .b(stage5_col99[4]),
        .s(ha_s5_c99_n22_s),
        .c_out(ha_s5_c99_n22_c)
    );

    ha ha_s5_c101_n23 (
        .a(stage5_col101[3]),
        .b(stage5_col101[4]),
        .s(ha_s5_c101_n23_s),
        .c_out(ha_s5_c101_n23_c)
    );

    ha ha_s5_c103_n24 (
        .a(stage5_col103[3]),
        .b(stage5_col103[4]),
        .s(ha_s5_c103_n24_s),
        .c_out(ha_s5_c103_n24_c)
    );

    ha ha_s5_c105_n25 (
        .a(stage5_col105[3]),
        .b(stage5_col105[4]),
        .s(ha_s5_c105_n25_s),
        .c_out(ha_s5_c105_n25_c)
    );

    ha ha_s5_c107_n26 (
        .a(stage5_col107[3]),
        .b(stage5_col107[4]),
        .s(ha_s5_c107_n26_s),
        .c_out(ha_s5_c107_n26_c)
    );

    ha ha_s5_c109_n27 (
        .a(stage5_col109[3]),
        .b(stage5_col109[4]),
        .s(ha_s5_c109_n27_s),
        .c_out(ha_s5_c109_n27_c)
    );

    ha ha_s5_c111_n28 (
        .a(stage5_col111[3]),
        .b(stage5_col111[4]),
        .s(ha_s5_c111_n28_s),
        .c_out(ha_s5_c111_n28_c)
    );

    ha ha_s5_c113_n29 (
        .a(stage5_col113[3]),
        .b(stage5_col113[4]),
        .s(ha_s5_c113_n29_s),
        .c_out(ha_s5_c113_n29_c)
    );

    ha ha_s5_c115_n30 (
        .a(stage5_col115[3]),
        .b(stage5_col115[4]),
        .s(ha_s5_c115_n30_s),
        .c_out(ha_s5_c115_n30_c)
    );

    ha ha_s5_c117_n31 (
        .a(stage5_col117[3]),
        .b(stage5_col117[4]),
        .s(ha_s5_c117_n31_s),
        .c_out(ha_s5_c117_n31_c)
    );

    ha ha_s5_c119_n32 (
        .a(stage5_col119[3]),
        .b(stage5_col119[4]),
        .s(ha_s5_c119_n32_s),
        .c_out(ha_s5_c119_n32_c)
    );

    ha ha_s5_c121_n33 (
        .a(stage5_col121[3]),
        .b(stage5_col121[4]),
        .s(ha_s5_c121_n33_s),
        .c_out(ha_s5_c121_n33_c)
    );

    ha ha_s5_c123_n34 (
        .a(stage5_col123[3]),
        .b(stage5_col123[4]),
        .s(ha_s5_c123_n34_s),
        .c_out(ha_s5_c123_n34_c)
    );

    ha ha_s5_c125_n35 (
        .a(stage5_col125[3]),
        .b(stage5_col125[4]),
        .s(ha_s5_c125_n35_s),
        .c_out(ha_s5_c125_n35_c)
    );

    // Map to Stage 6 columns
    generate
        if (PIPE) begin : gen_stage6_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage6_col0[0] <= 1'b0;
                    stage6_col1[0] <= 1'b0;
                    stage6_col2[0] <= 1'b0;
                    stage6_col3[0] <= 1'b0;
                    stage6_col4[0] <= 1'b0;
                    stage6_col5[0] <= 1'b0;
                    stage6_col6[0] <= 1'b0;
                    stage6_col6[1] <= 1'b0;
                    stage6_col7[0] <= 1'b0;
                    stage6_col8[0] <= 1'b0;
                    stage6_col8[1] <= 1'b0;
                    stage6_col8[2] <= 1'b0;
                    stage6_col9[0] <= 1'b0;
                    stage6_col9[1] <= 1'b0;
                    stage6_col10[0] <= 1'b0;
                    stage6_col10[1] <= 1'b0;
                    stage6_col11[0] <= 1'b0;
                    stage6_col11[1] <= 1'b0;
                    stage6_col12[0] <= 1'b0;
                    stage6_col12[1] <= 1'b0;
                    stage6_col13[0] <= 1'b0;
                    stage6_col13[1] <= 1'b0;
                    stage6_col14[0] <= 1'b0;
                    stage6_col14[1] <= 1'b0;
                    stage6_col15[0] <= 1'b0;
                    stage6_col15[1] <= 1'b0;
                    stage6_col16[0] <= 1'b0;
                    stage6_col16[1] <= 1'b0;
                    stage6_col17[0] <= 1'b0;
                    stage6_col17[1] <= 1'b0;
                    stage6_col18[0] <= 1'b0;
                    stage6_col18[1] <= 1'b0;
                    stage6_col19[0] <= 1'b0;
                    stage6_col19[1] <= 1'b0;
                    stage6_col20[0] <= 1'b0;
                    stage6_col20[1] <= 1'b0;
                    stage6_col21[0] <= 1'b0;
                    stage6_col21[1] <= 1'b0;
                    stage6_col22[0] <= 1'b0;
                    stage6_col22[1] <= 1'b0;
                    stage6_col23[0] <= 1'b0;
                    stage6_col23[1] <= 1'b0;
                    stage6_col24[0] <= 1'b0;
                    stage6_col24[1] <= 1'b0;
                    stage6_col25[0] <= 1'b0;
                    stage6_col25[1] <= 1'b0;
                    stage6_col26[0] <= 1'b0;
                    stage6_col26[1] <= 1'b0;
                    stage6_col27[0] <= 1'b0;
                    stage6_col27[1] <= 1'b0;
                    stage6_col28[0] <= 1'b0;
                    stage6_col28[1] <= 1'b0;
                    stage6_col29[0] <= 1'b0;
                    stage6_col29[1] <= 1'b0;
                    stage6_col30[0] <= 1'b0;
                    stage6_col30[1] <= 1'b0;
                    stage6_col31[0] <= 1'b0;
                    stage6_col31[1] <= 1'b0;
                    stage6_col32[0] <= 1'b0;
                    stage6_col32[1] <= 1'b0;
                    stage6_col33[0] <= 1'b0;
                    stage6_col33[1] <= 1'b0;
                    stage6_col34[0] <= 1'b0;
                    stage6_col34[1] <= 1'b0;
                    stage6_col35[0] <= 1'b0;
                    stage6_col35[1] <= 1'b0;
                    stage6_col36[0] <= 1'b0;
                    stage6_col36[1] <= 1'b0;
                    stage6_col37[0] <= 1'b0;
                    stage6_col37[1] <= 1'b0;
                    stage6_col38[0] <= 1'b0;
                    stage6_col38[1] <= 1'b0;
                    stage6_col39[0] <= 1'b0;
                    stage6_col39[1] <= 1'b0;
                    stage6_col40[0] <= 1'b0;
                    stage6_col40[1] <= 1'b0;
                    stage6_col41[0] <= 1'b0;
                    stage6_col41[1] <= 1'b0;
                    stage6_col41[2] <= 1'b0;
                    stage6_col41[3] <= 1'b0;
                    stage6_col42[0] <= 1'b0;
                    stage6_col42[1] <= 1'b0;
                    stage6_col42[2] <= 1'b0;
                    stage6_col43[0] <= 1'b0;
                    stage6_col43[1] <= 1'b0;
                    stage6_col43[2] <= 1'b0;
                    stage6_col44[0] <= 1'b0;
                    stage6_col44[1] <= 1'b0;
                    stage6_col44[2] <= 1'b0;
                    stage6_col45[0] <= 1'b0;
                    stage6_col45[1] <= 1'b0;
                    stage6_col45[2] <= 1'b0;
                    stage6_col46[0] <= 1'b0;
                    stage6_col46[1] <= 1'b0;
                    stage6_col46[2] <= 1'b0;
                    stage6_col47[0] <= 1'b0;
                    stage6_col47[1] <= 1'b0;
                    stage6_col47[2] <= 1'b0;
                    stage6_col48[0] <= 1'b0;
                    stage6_col48[1] <= 1'b0;
                    stage6_col48[2] <= 1'b0;
                    stage6_col49[0] <= 1'b0;
                    stage6_col49[1] <= 1'b0;
                    stage6_col49[2] <= 1'b0;
                    stage6_col50[0] <= 1'b0;
                    stage6_col50[1] <= 1'b0;
                    stage6_col50[2] <= 1'b0;
                    stage6_col51[0] <= 1'b0;
                    stage6_col51[1] <= 1'b0;
                    stage6_col51[2] <= 1'b0;
                    stage6_col52[0] <= 1'b0;
                    stage6_col52[1] <= 1'b0;
                    stage6_col52[2] <= 1'b0;
                    stage6_col53[0] <= 1'b0;
                    stage6_col53[1] <= 1'b0;
                    stage6_col53[2] <= 1'b0;
                    stage6_col54[0] <= 1'b0;
                    stage6_col54[1] <= 1'b0;
                    stage6_col54[2] <= 1'b0;
                    stage6_col55[0] <= 1'b0;
                    stage6_col55[1] <= 1'b0;
                    stage6_col55[2] <= 1'b0;
                    stage6_col56[0] <= 1'b0;
                    stage6_col56[1] <= 1'b0;
                    stage6_col56[2] <= 1'b0;
                    stage6_col57[0] <= 1'b0;
                    stage6_col57[1] <= 1'b0;
                    stage6_col57[2] <= 1'b0;
                    stage6_col58[0] <= 1'b0;
                    stage6_col58[1] <= 1'b0;
                    stage6_col58[2] <= 1'b0;
                    stage6_col59[0] <= 1'b0;
                    stage6_col59[1] <= 1'b0;
                    stage6_col59[2] <= 1'b0;
                    stage6_col60[0] <= 1'b0;
                    stage6_col60[1] <= 1'b0;
                    stage6_col60[2] <= 1'b0;
                    stage6_col60[3] <= 1'b0;
                    stage6_col61[0] <= 1'b0;
                    stage6_col61[1] <= 1'b0;
                    stage6_col61[2] <= 1'b0;
                    stage6_col61[3] <= 1'b0;
                    stage6_col62[0] <= 1'b0;
                    stage6_col62[1] <= 1'b0;
                    stage6_col62[2] <= 1'b0;
                    stage6_col62[3] <= 1'b0;
                    stage6_col63[0] <= 1'b0;
                    stage6_col63[1] <= 1'b0;
                    stage6_col63[2] <= 1'b0;
                    stage6_col63[3] <= 1'b0;
                    stage6_col64[0] <= 1'b0;
                    stage6_col64[1] <= 1'b0;
                    stage6_col64[2] <= 1'b0;
                    stage6_col64[3] <= 1'b0;
                    stage6_col65[0] <= 1'b0;
                    stage6_col65[1] <= 1'b0;
                    stage6_col65[2] <= 1'b0;
                    stage6_col65[3] <= 1'b0;
                    stage6_col66[0] <= 1'b0;
                    stage6_col66[1] <= 1'b0;
                    stage6_col66[2] <= 1'b0;
                    stage6_col66[3] <= 1'b0;
                    stage6_col67[0] <= 1'b0;
                    stage6_col67[1] <= 1'b0;
                    stage6_col67[2] <= 1'b0;
                    stage6_col67[3] <= 1'b0;
                    stage6_col68[0] <= 1'b0;
                    stage6_col68[1] <= 1'b0;
                    stage6_col68[2] <= 1'b0;
                    stage6_col68[3] <= 1'b0;
                    stage6_col69[0] <= 1'b0;
                    stage6_col69[1] <= 1'b0;
                    stage6_col69[2] <= 1'b0;
                    stage6_col69[3] <= 1'b0;
                    stage6_col70[0] <= 1'b0;
                    stage6_col70[1] <= 1'b0;
                    stage6_col70[2] <= 1'b0;
                    stage6_col70[3] <= 1'b0;
                    stage6_col71[0] <= 1'b0;
                    stage6_col71[1] <= 1'b0;
                    stage6_col71[2] <= 1'b0;
                    stage6_col71[3] <= 1'b0;
                    stage6_col72[0] <= 1'b0;
                    stage6_col72[1] <= 1'b0;
                    stage6_col72[2] <= 1'b0;
                    stage6_col72[3] <= 1'b0;
                    stage6_col73[0] <= 1'b0;
                    stage6_col73[1] <= 1'b0;
                    stage6_col73[2] <= 1'b0;
                    stage6_col73[3] <= 1'b0;
                    stage6_col74[0] <= 1'b0;
                    stage6_col74[1] <= 1'b0;
                    stage6_col74[2] <= 1'b0;
                    stage6_col74[3] <= 1'b0;
                    stage6_col75[0] <= 1'b0;
                    stage6_col75[1] <= 1'b0;
                    stage6_col75[2] <= 1'b0;
                    stage6_col75[3] <= 1'b0;
                    stage6_col76[0] <= 1'b0;
                    stage6_col76[1] <= 1'b0;
                    stage6_col76[2] <= 1'b0;
                    stage6_col76[3] <= 1'b0;
                    stage6_col77[0] <= 1'b0;
                    stage6_col77[1] <= 1'b0;
                    stage6_col77[2] <= 1'b0;
                    stage6_col77[3] <= 1'b0;
                    stage6_col78[0] <= 1'b0;
                    stage6_col78[1] <= 1'b0;
                    stage6_col78[2] <= 1'b0;
                    stage6_col78[3] <= 1'b0;
                    stage6_col79[0] <= 1'b0;
                    stage6_col79[1] <= 1'b0;
                    stage6_col79[2] <= 1'b0;
                    stage6_col79[3] <= 1'b0;
                    stage6_col80[0] <= 1'b0;
                    stage6_col80[1] <= 1'b0;
                    stage6_col80[2] <= 1'b0;
                    stage6_col80[3] <= 1'b0;
                    stage6_col81[0] <= 1'b0;
                    stage6_col81[1] <= 1'b0;
                    stage6_col81[2] <= 1'b0;
                    stage6_col81[3] <= 1'b0;
                    stage6_col82[0] <= 1'b0;
                    stage6_col82[1] <= 1'b0;
                    stage6_col82[2] <= 1'b0;
                    stage6_col82[3] <= 1'b0;
                    stage6_col83[0] <= 1'b0;
                    stage6_col83[1] <= 1'b0;
                    stage6_col83[2] <= 1'b0;
                    stage6_col83[3] <= 1'b0;
                    stage6_col84[0] <= 1'b0;
                    stage6_col84[1] <= 1'b0;
                    stage6_col84[2] <= 1'b0;
                    stage6_col84[3] <= 1'b0;
                    stage6_col85[0] <= 1'b0;
                    stage6_col85[1] <= 1'b0;
                    stage6_col85[2] <= 1'b0;
                    stage6_col85[3] <= 1'b0;
                    stage6_col86[0] <= 1'b0;
                    stage6_col86[1] <= 1'b0;
                    stage6_col86[2] <= 1'b0;
                    stage6_col86[3] <= 1'b0;
                    stage6_col87[0] <= 1'b0;
                    stage6_col87[1] <= 1'b0;
                    stage6_col87[2] <= 1'b0;
                    stage6_col87[3] <= 1'b0;
                    stage6_col88[0] <= 1'b0;
                    stage6_col88[1] <= 1'b0;
                    stage6_col88[2] <= 1'b0;
                    stage6_col88[3] <= 1'b0;
                    stage6_col89[0] <= 1'b0;
                    stage6_col89[1] <= 1'b0;
                    stage6_col89[2] <= 1'b0;
                    stage6_col89[3] <= 1'b0;
                    stage6_col90[0] <= 1'b0;
                    stage6_col90[1] <= 1'b0;
                    stage6_col90[2] <= 1'b0;
                    stage6_col90[3] <= 1'b0;
                    stage6_col91[0] <= 1'b0;
                    stage6_col91[1] <= 1'b0;
                    stage6_col91[2] <= 1'b0;
                    stage6_col91[3] <= 1'b0;
                    stage6_col92[0] <= 1'b0;
                    stage6_col92[1] <= 1'b0;
                    stage6_col92[2] <= 1'b0;
                    stage6_col92[3] <= 1'b0;
                    stage6_col93[0] <= 1'b0;
                    stage6_col93[1] <= 1'b0;
                    stage6_col93[2] <= 1'b0;
                    stage6_col93[3] <= 1'b0;
                    stage6_col94[0] <= 1'b0;
                    stage6_col94[1] <= 1'b0;
                    stage6_col94[2] <= 1'b0;
                    stage6_col94[3] <= 1'b0;
                    stage6_col95[0] <= 1'b0;
                    stage6_col95[1] <= 1'b0;
                    stage6_col95[2] <= 1'b0;
                    stage6_col95[3] <= 1'b0;
                    stage6_col96[0] <= 1'b0;
                    stage6_col96[1] <= 1'b0;
                    stage6_col96[2] <= 1'b0;
                    stage6_col96[3] <= 1'b0;
                    stage6_col97[0] <= 1'b0;
                    stage6_col97[1] <= 1'b0;
                    stage6_col97[2] <= 1'b0;
                    stage6_col97[3] <= 1'b0;
                    stage6_col98[0] <= 1'b0;
                    stage6_col98[1] <= 1'b0;
                    stage6_col98[2] <= 1'b0;
                    stage6_col98[3] <= 1'b0;
                    stage6_col99[0] <= 1'b0;
                    stage6_col99[1] <= 1'b0;
                    stage6_col99[2] <= 1'b0;
                    stage6_col99[3] <= 1'b0;
                    stage6_col100[0] <= 1'b0;
                    stage6_col100[1] <= 1'b0;
                    stage6_col100[2] <= 1'b0;
                    stage6_col100[3] <= 1'b0;
                    stage6_col101[0] <= 1'b0;
                    stage6_col101[1] <= 1'b0;
                    stage6_col101[2] <= 1'b0;
                    stage6_col101[3] <= 1'b0;
                    stage6_col102[0] <= 1'b0;
                    stage6_col102[1] <= 1'b0;
                    stage6_col102[2] <= 1'b0;
                    stage6_col102[3] <= 1'b0;
                    stage6_col103[0] <= 1'b0;
                    stage6_col103[1] <= 1'b0;
                    stage6_col103[2] <= 1'b0;
                    stage6_col103[3] <= 1'b0;
                    stage6_col104[0] <= 1'b0;
                    stage6_col104[1] <= 1'b0;
                    stage6_col104[2] <= 1'b0;
                    stage6_col104[3] <= 1'b0;
                    stage6_col105[0] <= 1'b0;
                    stage6_col105[1] <= 1'b0;
                    stage6_col105[2] <= 1'b0;
                    stage6_col105[3] <= 1'b0;
                    stage6_col106[0] <= 1'b0;
                    stage6_col106[1] <= 1'b0;
                    stage6_col106[2] <= 1'b0;
                    stage6_col106[3] <= 1'b0;
                    stage6_col107[0] <= 1'b0;
                    stage6_col107[1] <= 1'b0;
                    stage6_col107[2] <= 1'b0;
                    stage6_col107[3] <= 1'b0;
                    stage6_col108[0] <= 1'b0;
                    stage6_col108[1] <= 1'b0;
                    stage6_col108[2] <= 1'b0;
                    stage6_col108[3] <= 1'b0;
                    stage6_col109[0] <= 1'b0;
                    stage6_col109[1] <= 1'b0;
                    stage6_col109[2] <= 1'b0;
                    stage6_col109[3] <= 1'b0;
                    stage6_col110[0] <= 1'b0;
                    stage6_col110[1] <= 1'b0;
                    stage6_col110[2] <= 1'b0;
                    stage6_col110[3] <= 1'b0;
                    stage6_col111[0] <= 1'b0;
                    stage6_col111[1] <= 1'b0;
                    stage6_col111[2] <= 1'b0;
                    stage6_col111[3] <= 1'b0;
                    stage6_col112[0] <= 1'b0;
                    stage6_col112[1] <= 1'b0;
                    stage6_col112[2] <= 1'b0;
                    stage6_col112[3] <= 1'b0;
                    stage6_col113[0] <= 1'b0;
                    stage6_col113[1] <= 1'b0;
                    stage6_col113[2] <= 1'b0;
                    stage6_col113[3] <= 1'b0;
                    stage6_col114[0] <= 1'b0;
                    stage6_col114[1] <= 1'b0;
                    stage6_col114[2] <= 1'b0;
                    stage6_col114[3] <= 1'b0;
                    stage6_col115[0] <= 1'b0;
                    stage6_col115[1] <= 1'b0;
                    stage6_col115[2] <= 1'b0;
                    stage6_col115[3] <= 1'b0;
                    stage6_col116[0] <= 1'b0;
                    stage6_col116[1] <= 1'b0;
                    stage6_col116[2] <= 1'b0;
                    stage6_col116[3] <= 1'b0;
                    stage6_col117[0] <= 1'b0;
                    stage6_col117[1] <= 1'b0;
                    stage6_col117[2] <= 1'b0;
                    stage6_col117[3] <= 1'b0;
                    stage6_col118[0] <= 1'b0;
                    stage6_col118[1] <= 1'b0;
                    stage6_col118[2] <= 1'b0;
                    stage6_col118[3] <= 1'b0;
                    stage6_col119[0] <= 1'b0;
                    stage6_col119[1] <= 1'b0;
                    stage6_col119[2] <= 1'b0;
                    stage6_col119[3] <= 1'b0;
                    stage6_col120[0] <= 1'b0;
                    stage6_col120[1] <= 1'b0;
                    stage6_col120[2] <= 1'b0;
                    stage6_col120[3] <= 1'b0;
                    stage6_col121[0] <= 1'b0;
                    stage6_col121[1] <= 1'b0;
                    stage6_col121[2] <= 1'b0;
                    stage6_col121[3] <= 1'b0;
                    stage6_col122[0] <= 1'b0;
                    stage6_col122[1] <= 1'b0;
                    stage6_col122[2] <= 1'b0;
                    stage6_col122[3] <= 1'b0;
                    stage6_col123[0] <= 1'b0;
                    stage6_col123[1] <= 1'b0;
                    stage6_col123[2] <= 1'b0;
                    stage6_col123[3] <= 1'b0;
                    stage6_col124[0] <= 1'b0;
                    stage6_col124[1] <= 1'b0;
                    stage6_col124[2] <= 1'b0;
                    stage6_col124[3] <= 1'b0;
                    stage6_col125[0] <= 1'b0;
                    stage6_col125[1] <= 1'b0;
                    stage6_col125[2] <= 1'b0;
                    stage6_col125[3] <= 1'b0;
                    stage6_col126[0] <= 1'b0;
                    stage6_col126[1] <= 1'b0;
                    stage6_col126[2] <= 1'b0;
                    stage6_col126[3] <= 1'b0;
                    stage6_col127[0] <= 1'b0;
                    stage6_col127[1] <= 1'b0;
                    stage6_col127[2] <= 1'b0;
                    stage6_col127[3] <= 1'b0;
                    stage6_col127[4] <= 1'b0;
                    stage6_col127[5] <= 1'b0;
                    stage6_col127[6] <= 1'b0;
                    stage6_col127[7] <= 1'b0;
                    stage6_col127[8] <= 1'b0;
                    stage6_col127[9] <= 1'b0;
                    stage6_col127[10] <= 1'b0;
                    stage6_col127[11] <= 1'b0;
                    stage6_col127[12] <= 1'b0;
                    stage6_col127[13] <= 1'b0;
                    stage6_col127[14] <= 1'b0;
                    stage6_col127[15] <= 1'b0;
                    stage6_col127[16] <= 1'b0;
                    stage6_col127[17] <= 1'b0;
                    stage6_col127[18] <= 1'b0;
                    stage6_col127[19] <= 1'b0;
                    stage6_col127[20] <= 1'b0;
                    stage6_col127[21] <= 1'b0;
                    stage6_col127[22] <= 1'b0;
                    stage6_col127[23] <= 1'b0;
                    stage6_col127[24] <= 1'b0;
                    stage6_col127[25] <= 1'b0;
                    stage6_col127[26] <= 1'b0;
                    stage6_col127[27] <= 1'b0;
                    stage6_col127[28] <= 1'b0;
                    stage6_col127[29] <= 1'b0;
                    stage6_col127[30] <= 1'b0;
                    stage6_col127[31] <= 1'b0;
                    stage6_col127[32] <= 1'b0;
                    stage6_col127[33] <= 1'b0;
                    stage6_col127[34] <= 1'b0;
                    stage6_col127[35] <= 1'b0;
                    stage6_col127[36] <= 1'b0;
                    stage6_col127[37] <= 1'b0;
                    stage6_col127[38] <= 1'b0;
                    stage6_col127[39] <= 1'b0;
                    stage6_col127[40] <= 1'b0;
                    stage6_col127[41] <= 1'b0;
                    stage6_col127[42] <= 1'b0;
                    stage6_col127[43] <= 1'b0;
                    stage6_col127[44] <= 1'b0;
                    stage6_col127[45] <= 1'b0;
                    stage6_col127[46] <= 1'b0;
                    stage6_col127[47] <= 1'b0;
                    stage6_col127[48] <= 1'b0;
                    stage6_col127[49] <= 1'b0;
                    stage6_col127[50] <= 1'b0;
                    stage6_col127[51] <= 1'b0;
                    stage6_col127[52] <= 1'b0;
                    stage6_col127[53] <= 1'b0;
                    stage6_col127[54] <= 1'b0;
                    stage6_col127[55] <= 1'b0;
                    stage6_col127[56] <= 1'b0;
                    stage6_col127[57] <= 1'b0;
                    stage6_col127[58] <= 1'b0;
                    stage6_col127[59] <= 1'b0;
                    stage6_col127[60] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage6_col0[0] <= stage5_col0[0];
                    stage6_col1[0] <= stage5_col1[0];
                    stage6_col2[0] <= stage5_col2[0];
                    stage6_col3[0] <= stage5_col3[0];
                    stage6_col4[0] <= stage5_col4[0];
                    stage6_col5[0] <= ha_s5_c5_n0_s;
                    stage6_col6[0] <= ha_s5_c5_n0_c;
                    stage6_col6[1] <= stage5_col6[0];
                    stage6_col7[0] <= fa_s5_c7_n0_s;
                    stage6_col8[0] <= fa_s5_c7_n0_c;
                    stage6_col8[1] <= stage5_col8[0];
                    stage6_col8[2] <= stage5_col8[1];
                    stage6_col9[0] <= stage5_col9[0];
                    stage6_col9[1] <= stage5_col9[1];
                    stage6_col10[0] <= stage5_col10[0];
                    stage6_col10[1] <= stage5_col10[1];
                    stage6_col11[0] <= stage5_col11[0];
                    stage6_col11[1] <= stage5_col11[1];
                    stage6_col12[0] <= stage5_col12[0];
                    stage6_col12[1] <= stage5_col12[1];
                    stage6_col13[0] <= stage5_col13[0];
                    stage6_col13[1] <= stage5_col13[1];
                    stage6_col14[0] <= stage5_col14[0];
                    stage6_col14[1] <= stage5_col14[1];
                    stage6_col15[0] <= stage5_col15[0];
                    stage6_col15[1] <= stage5_col15[1];
                    stage6_col16[0] <= stage5_col16[0];
                    stage6_col16[1] <= stage5_col16[1];
                    stage6_col17[0] <= stage5_col17[0];
                    stage6_col17[1] <= stage5_col17[1];
                    stage6_col18[0] <= stage5_col18[0];
                    stage6_col18[1] <= stage5_col18[1];
                    stage6_col19[0] <= stage5_col19[0];
                    stage6_col19[1] <= stage5_col19[1];
                    stage6_col20[0] <= stage5_col20[0];
                    stage6_col20[1] <= stage5_col20[1];
                    stage6_col21[0] <= stage5_col21[0];
                    stage6_col21[1] <= stage5_col21[1];
                    stage6_col22[0] <= stage5_col22[0];
                    stage6_col22[1] <= stage5_col22[1];
                    stage6_col23[0] <= stage5_col23[0];
                    stage6_col23[1] <= stage5_col23[1];
                    stage6_col24[0] <= stage5_col24[0];
                    stage6_col24[1] <= stage5_col24[1];
                    stage6_col25[0] <= stage5_col25[0];
                    stage6_col25[1] <= stage5_col25[1];
                    stage6_col26[0] <= stage5_col26[0];
                    stage6_col26[1] <= stage5_col26[1];
                    stage6_col27[0] <= stage5_col27[0];
                    stage6_col27[1] <= stage5_col27[1];
                    stage6_col28[0] <= fa_s5_c28_n1_s;
                    stage6_col28[1] <= stage5_col28[3];
                    stage6_col29[0] <= fa_s5_c28_n1_c;
                    stage6_col29[1] <= fa_s5_c29_n2_s;
                    stage6_col30[0] <= fa_s5_c29_n2_c;
                    stage6_col30[1] <= fa_s5_c30_n3_s;
                    stage6_col31[0] <= fa_s5_c30_n3_c;
                    stage6_col31[1] <= fa_s5_c31_n4_s;
                    stage6_col32[0] <= fa_s5_c31_n4_c;
                    stage6_col32[1] <= fa_s5_c32_n5_s;
                    stage6_col33[0] <= fa_s5_c32_n5_c;
                    stage6_col33[1] <= fa_s5_c33_n6_s;
                    stage6_col34[0] <= fa_s5_c33_n6_c;
                    stage6_col34[1] <= fa_s5_c34_n7_s;
                    stage6_col35[0] <= fa_s5_c34_n7_c;
                    stage6_col35[1] <= fa_s5_c35_n8_s;
                    stage6_col36[0] <= fa_s5_c35_n8_c;
                    stage6_col36[1] <= fa_s5_c36_n9_s;
                    stage6_col37[0] <= fa_s5_c36_n9_c;
                    stage6_col37[1] <= fa_s5_c37_n10_s;
                    stage6_col38[0] <= fa_s5_c37_n10_c;
                    stage6_col38[1] <= fa_s5_c38_n11_s;
                    stage6_col39[0] <= fa_s5_c38_n11_c;
                    stage6_col39[1] <= fa_s5_c39_n12_s;
                    stage6_col40[0] <= fa_s5_c39_n12_c;
                    stage6_col40[1] <= fa_s5_c40_n13_s;
                    stage6_col41[0] <= fa_s5_c40_n13_c;
                    stage6_col41[1] <= fa_s5_c41_n14_s;
                    stage6_col41[2] <= stage5_col41[3];
                    stage6_col41[3] <= stage5_col41[4];
                    stage6_col42[0] <= fa_s5_c41_n14_c;
                    stage6_col42[1] <= fa_s5_c42_n15_s;
                    stage6_col42[2] <= stage5_col42[3];
                    stage6_col43[0] <= fa_s5_c42_n15_c;
                    stage6_col43[1] <= fa_s5_c43_n16_s;
                    stage6_col43[2] <= stage5_col43[3];
                    stage6_col44[0] <= fa_s5_c43_n16_c;
                    stage6_col44[1] <= fa_s5_c44_n17_s;
                    stage6_col44[2] <= stage5_col44[3];
                    stage6_col45[0] <= fa_s5_c44_n17_c;
                    stage6_col45[1] <= fa_s5_c45_n18_s;
                    stage6_col45[2] <= stage5_col45[3];
                    stage6_col46[0] <= fa_s5_c45_n18_c;
                    stage6_col46[1] <= fa_s5_c46_n19_s;
                    stage6_col46[2] <= stage5_col46[3];
                    stage6_col47[0] <= fa_s5_c46_n19_c;
                    stage6_col47[1] <= fa_s5_c47_n20_s;
                    stage6_col47[2] <= stage5_col47[3];
                    stage6_col48[0] <= fa_s5_c47_n20_c;
                    stage6_col48[1] <= fa_s5_c48_n21_s;
                    stage6_col48[2] <= stage5_col48[3];
                    stage6_col49[0] <= fa_s5_c48_n21_c;
                    stage6_col49[1] <= fa_s5_c49_n22_s;
                    stage6_col49[2] <= stage5_col49[3];
                    stage6_col50[0] <= fa_s5_c49_n22_c;
                    stage6_col50[1] <= fa_s5_c50_n23_s;
                    stage6_col50[2] <= stage5_col50[3];
                    stage6_col51[0] <= fa_s5_c50_n23_c;
                    stage6_col51[1] <= fa_s5_c51_n24_s;
                    stage6_col51[2] <= stage5_col51[3];
                    stage6_col52[0] <= fa_s5_c51_n24_c;
                    stage6_col52[1] <= fa_s5_c52_n25_s;
                    stage6_col52[2] <= stage5_col52[3];
                    stage6_col53[0] <= fa_s5_c52_n25_c;
                    stage6_col53[1] <= fa_s5_c53_n26_s;
                    stage6_col53[2] <= stage5_col53[3];
                    stage6_col54[0] <= fa_s5_c53_n26_c;
                    stage6_col54[1] <= fa_s5_c54_n27_s;
                    stage6_col54[2] <= stage5_col54[3];
                    stage6_col55[0] <= fa_s5_c54_n27_c;
                    stage6_col55[1] <= fa_s5_c55_n28_s;
                    stage6_col55[2] <= stage5_col55[3];
                    stage6_col56[0] <= fa_s5_c55_n28_c;
                    stage6_col56[1] <= fa_s5_c56_n29_s;
                    stage6_col56[2] <= stage5_col56[3];
                    stage6_col57[0] <= fa_s5_c56_n29_c;
                    stage6_col57[1] <= fa_s5_c57_n30_s;
                    stage6_col57[2] <= stage5_col57[3];
                    stage6_col58[0] <= fa_s5_c57_n30_c;
                    stage6_col58[1] <= fa_s5_c58_n31_s;
                    stage6_col58[2] <= stage5_col58[3];
                    stage6_col59[0] <= fa_s5_c58_n31_c;
                    stage6_col59[1] <= fa_s5_c59_n32_s;
                    stage6_col59[2] <= fa_s5_c59_n33_s;
                    stage6_col60[0] <= fa_s5_c59_n32_c;
                    stage6_col60[1] <= fa_s5_c59_n33_c;
                    stage6_col60[2] <= fa_s5_c60_n34_s;
                    stage6_col60[3] <= ha_s5_c60_n1_s;
                    stage6_col61[0] <= fa_s5_c60_n34_c;
                    stage6_col61[1] <= ha_s5_c60_n1_c;
                    stage6_col61[2] <= fa_s5_c61_n35_s;
                    stage6_col61[3] <= ha_s5_c61_n2_s;
                    stage6_col62[0] <= fa_s5_c61_n35_c;
                    stage6_col62[1] <= ha_s5_c61_n2_c;
                    stage6_col62[2] <= fa_s5_c62_n36_s;
                    stage6_col62[3] <= ha_s5_c62_n3_s;
                    stage6_col63[0] <= fa_s5_c62_n36_c;
                    stage6_col63[1] <= ha_s5_c62_n3_c;
                    stage6_col63[2] <= fa_s5_c63_n37_s;
                    stage6_col63[3] <= ha_s5_c63_n4_s;
                    stage6_col64[0] <= fa_s5_c63_n37_c;
                    stage6_col64[1] <= ha_s5_c63_n4_c;
                    stage6_col64[2] <= fa_s5_c64_n38_s;
                    stage6_col64[3] <= fa_s5_c64_n39_s;
                    stage6_col65[0] <= fa_s5_c64_n38_c;
                    stage6_col65[1] <= fa_s5_c64_n39_c;
                    stage6_col65[2] <= fa_s5_c65_n40_s;
                    stage6_col65[3] <= ha_s5_c65_n5_s;
                    stage6_col66[0] <= fa_s5_c65_n40_c;
                    stage6_col66[1] <= ha_s5_c65_n5_c;
                    stage6_col66[2] <= fa_s5_c66_n41_s;
                    stage6_col66[3] <= fa_s5_c66_n42_s;
                    stage6_col67[0] <= fa_s5_c66_n41_c;
                    stage6_col67[1] <= fa_s5_c66_n42_c;
                    stage6_col67[2] <= fa_s5_c67_n43_s;
                    stage6_col67[3] <= ha_s5_c67_n6_s;
                    stage6_col68[0] <= fa_s5_c67_n43_c;
                    stage6_col68[1] <= ha_s5_c67_n6_c;
                    stage6_col68[2] <= fa_s5_c68_n44_s;
                    stage6_col68[3] <= fa_s5_c68_n45_s;
                    stage6_col69[0] <= fa_s5_c68_n44_c;
                    stage6_col69[1] <= fa_s5_c68_n45_c;
                    stage6_col69[2] <= fa_s5_c69_n46_s;
                    stage6_col69[3] <= ha_s5_c69_n7_s;
                    stage6_col70[0] <= fa_s5_c69_n46_c;
                    stage6_col70[1] <= ha_s5_c69_n7_c;
                    stage6_col70[2] <= fa_s5_c70_n47_s;
                    stage6_col70[3] <= fa_s5_c70_n48_s;
                    stage6_col71[0] <= fa_s5_c70_n47_c;
                    stage6_col71[1] <= fa_s5_c70_n48_c;
                    stage6_col71[2] <= fa_s5_c71_n49_s;
                    stage6_col71[3] <= ha_s5_c71_n8_s;
                    stage6_col72[0] <= fa_s5_c71_n49_c;
                    stage6_col72[1] <= ha_s5_c71_n8_c;
                    stage6_col72[2] <= fa_s5_c72_n50_s;
                    stage6_col72[3] <= fa_s5_c72_n51_s;
                    stage6_col73[0] <= fa_s5_c72_n50_c;
                    stage6_col73[1] <= fa_s5_c72_n51_c;
                    stage6_col73[2] <= fa_s5_c73_n52_s;
                    stage6_col73[3] <= ha_s5_c73_n9_s;
                    stage6_col74[0] <= fa_s5_c73_n52_c;
                    stage6_col74[1] <= ha_s5_c73_n9_c;
                    stage6_col74[2] <= fa_s5_c74_n53_s;
                    stage6_col74[3] <= fa_s5_c74_n54_s;
                    stage6_col75[0] <= fa_s5_c74_n53_c;
                    stage6_col75[1] <= fa_s5_c74_n54_c;
                    stage6_col75[2] <= fa_s5_c75_n55_s;
                    stage6_col75[3] <= ha_s5_c75_n10_s;
                    stage6_col76[0] <= fa_s5_c75_n55_c;
                    stage6_col76[1] <= ha_s5_c75_n10_c;
                    stage6_col76[2] <= fa_s5_c76_n56_s;
                    stage6_col76[3] <= fa_s5_c76_n57_s;
                    stage6_col77[0] <= fa_s5_c76_n56_c;
                    stage6_col77[1] <= fa_s5_c76_n57_c;
                    stage6_col77[2] <= fa_s5_c77_n58_s;
                    stage6_col77[3] <= ha_s5_c77_n11_s;
                    stage6_col78[0] <= fa_s5_c77_n58_c;
                    stage6_col78[1] <= ha_s5_c77_n11_c;
                    stage6_col78[2] <= fa_s5_c78_n59_s;
                    stage6_col78[3] <= fa_s5_c78_n60_s;
                    stage6_col79[0] <= fa_s5_c78_n59_c;
                    stage6_col79[1] <= fa_s5_c78_n60_c;
                    stage6_col79[2] <= fa_s5_c79_n61_s;
                    stage6_col79[3] <= ha_s5_c79_n12_s;
                    stage6_col80[0] <= fa_s5_c79_n61_c;
                    stage6_col80[1] <= ha_s5_c79_n12_c;
                    stage6_col80[2] <= fa_s5_c80_n62_s;
                    stage6_col80[3] <= fa_s5_c80_n63_s;
                    stage6_col81[0] <= fa_s5_c80_n62_c;
                    stage6_col81[1] <= fa_s5_c80_n63_c;
                    stage6_col81[2] <= fa_s5_c81_n64_s;
                    stage6_col81[3] <= ha_s5_c81_n13_s;
                    stage6_col82[0] <= fa_s5_c81_n64_c;
                    stage6_col82[1] <= ha_s5_c81_n13_c;
                    stage6_col82[2] <= fa_s5_c82_n65_s;
                    stage6_col82[3] <= fa_s5_c82_n66_s;
                    stage6_col83[0] <= fa_s5_c82_n65_c;
                    stage6_col83[1] <= fa_s5_c82_n66_c;
                    stage6_col83[2] <= fa_s5_c83_n67_s;
                    stage6_col83[3] <= ha_s5_c83_n14_s;
                    stage6_col84[0] <= fa_s5_c83_n67_c;
                    stage6_col84[1] <= ha_s5_c83_n14_c;
                    stage6_col84[2] <= fa_s5_c84_n68_s;
                    stage6_col84[3] <= fa_s5_c84_n69_s;
                    stage6_col85[0] <= fa_s5_c84_n68_c;
                    stage6_col85[1] <= fa_s5_c84_n69_c;
                    stage6_col85[2] <= fa_s5_c85_n70_s;
                    stage6_col85[3] <= ha_s5_c85_n15_s;
                    stage6_col86[0] <= fa_s5_c85_n70_c;
                    stage6_col86[1] <= ha_s5_c85_n15_c;
                    stage6_col86[2] <= fa_s5_c86_n71_s;
                    stage6_col86[3] <= fa_s5_c86_n72_s;
                    stage6_col87[0] <= fa_s5_c86_n71_c;
                    stage6_col87[1] <= fa_s5_c86_n72_c;
                    stage6_col87[2] <= fa_s5_c87_n73_s;
                    stage6_col87[3] <= ha_s5_c87_n16_s;
                    stage6_col88[0] <= fa_s5_c87_n73_c;
                    stage6_col88[1] <= ha_s5_c87_n16_c;
                    stage6_col88[2] <= fa_s5_c88_n74_s;
                    stage6_col88[3] <= fa_s5_c88_n75_s;
                    stage6_col89[0] <= fa_s5_c88_n74_c;
                    stage6_col89[1] <= fa_s5_c88_n75_c;
                    stage6_col89[2] <= fa_s5_c89_n76_s;
                    stage6_col89[3] <= ha_s5_c89_n17_s;
                    stage6_col90[0] <= fa_s5_c89_n76_c;
                    stage6_col90[1] <= ha_s5_c89_n17_c;
                    stage6_col90[2] <= fa_s5_c90_n77_s;
                    stage6_col90[3] <= fa_s5_c90_n78_s;
                    stage6_col91[0] <= fa_s5_c90_n77_c;
                    stage6_col91[1] <= fa_s5_c90_n78_c;
                    stage6_col91[2] <= fa_s5_c91_n79_s;
                    stage6_col91[3] <= ha_s5_c91_n18_s;
                    stage6_col92[0] <= fa_s5_c91_n79_c;
                    stage6_col92[1] <= ha_s5_c91_n18_c;
                    stage6_col92[2] <= fa_s5_c92_n80_s;
                    stage6_col92[3] <= fa_s5_c92_n81_s;
                    stage6_col93[0] <= fa_s5_c92_n80_c;
                    stage6_col93[1] <= fa_s5_c92_n81_c;
                    stage6_col93[2] <= fa_s5_c93_n82_s;
                    stage6_col93[3] <= ha_s5_c93_n19_s;
                    stage6_col94[0] <= fa_s5_c93_n82_c;
                    stage6_col94[1] <= ha_s5_c93_n19_c;
                    stage6_col94[2] <= fa_s5_c94_n83_s;
                    stage6_col94[3] <= fa_s5_c94_n84_s;
                    stage6_col95[0] <= fa_s5_c94_n83_c;
                    stage6_col95[1] <= fa_s5_c94_n84_c;
                    stage6_col95[2] <= fa_s5_c95_n85_s;
                    stage6_col95[3] <= ha_s5_c95_n20_s;
                    stage6_col96[0] <= fa_s5_c95_n85_c;
                    stage6_col96[1] <= ha_s5_c95_n20_c;
                    stage6_col96[2] <= fa_s5_c96_n86_s;
                    stage6_col96[3] <= fa_s5_c96_n87_s;
                    stage6_col97[0] <= fa_s5_c96_n86_c;
                    stage6_col97[1] <= fa_s5_c96_n87_c;
                    stage6_col97[2] <= fa_s5_c97_n88_s;
                    stage6_col97[3] <= ha_s5_c97_n21_s;
                    stage6_col98[0] <= fa_s5_c97_n88_c;
                    stage6_col98[1] <= ha_s5_c97_n21_c;
                    stage6_col98[2] <= fa_s5_c98_n89_s;
                    stage6_col98[3] <= fa_s5_c98_n90_s;
                    stage6_col99[0] <= fa_s5_c98_n89_c;
                    stage6_col99[1] <= fa_s5_c98_n90_c;
                    stage6_col99[2] <= fa_s5_c99_n91_s;
                    stage6_col99[3] <= ha_s5_c99_n22_s;
                    stage6_col100[0] <= fa_s5_c99_n91_c;
                    stage6_col100[1] <= ha_s5_c99_n22_c;
                    stage6_col100[2] <= fa_s5_c100_n92_s;
                    stage6_col100[3] <= fa_s5_c100_n93_s;
                    stage6_col101[0] <= fa_s5_c100_n92_c;
                    stage6_col101[1] <= fa_s5_c100_n93_c;
                    stage6_col101[2] <= fa_s5_c101_n94_s;
                    stage6_col101[3] <= ha_s5_c101_n23_s;
                    stage6_col102[0] <= fa_s5_c101_n94_c;
                    stage6_col102[1] <= ha_s5_c101_n23_c;
                    stage6_col102[2] <= fa_s5_c102_n95_s;
                    stage6_col102[3] <= fa_s5_c102_n96_s;
                    stage6_col103[0] <= fa_s5_c102_n95_c;
                    stage6_col103[1] <= fa_s5_c102_n96_c;
                    stage6_col103[2] <= fa_s5_c103_n97_s;
                    stage6_col103[3] <= ha_s5_c103_n24_s;
                    stage6_col104[0] <= fa_s5_c103_n97_c;
                    stage6_col104[1] <= ha_s5_c103_n24_c;
                    stage6_col104[2] <= fa_s5_c104_n98_s;
                    stage6_col104[3] <= fa_s5_c104_n99_s;
                    stage6_col105[0] <= fa_s5_c104_n98_c;
                    stage6_col105[1] <= fa_s5_c104_n99_c;
                    stage6_col105[2] <= fa_s5_c105_n100_s;
                    stage6_col105[3] <= ha_s5_c105_n25_s;
                    stage6_col106[0] <= fa_s5_c105_n100_c;
                    stage6_col106[1] <= ha_s5_c105_n25_c;
                    stage6_col106[2] <= fa_s5_c106_n101_s;
                    stage6_col106[3] <= fa_s5_c106_n102_s;
                    stage6_col107[0] <= fa_s5_c106_n101_c;
                    stage6_col107[1] <= fa_s5_c106_n102_c;
                    stage6_col107[2] <= fa_s5_c107_n103_s;
                    stage6_col107[3] <= ha_s5_c107_n26_s;
                    stage6_col108[0] <= fa_s5_c107_n103_c;
                    stage6_col108[1] <= ha_s5_c107_n26_c;
                    stage6_col108[2] <= fa_s5_c108_n104_s;
                    stage6_col108[3] <= fa_s5_c108_n105_s;
                    stage6_col109[0] <= fa_s5_c108_n104_c;
                    stage6_col109[1] <= fa_s5_c108_n105_c;
                    stage6_col109[2] <= fa_s5_c109_n106_s;
                    stage6_col109[3] <= ha_s5_c109_n27_s;
                    stage6_col110[0] <= fa_s5_c109_n106_c;
                    stage6_col110[1] <= ha_s5_c109_n27_c;
                    stage6_col110[2] <= fa_s5_c110_n107_s;
                    stage6_col110[3] <= fa_s5_c110_n108_s;
                    stage6_col111[0] <= fa_s5_c110_n107_c;
                    stage6_col111[1] <= fa_s5_c110_n108_c;
                    stage6_col111[2] <= fa_s5_c111_n109_s;
                    stage6_col111[3] <= ha_s5_c111_n28_s;
                    stage6_col112[0] <= fa_s5_c111_n109_c;
                    stage6_col112[1] <= ha_s5_c111_n28_c;
                    stage6_col112[2] <= fa_s5_c112_n110_s;
                    stage6_col112[3] <= fa_s5_c112_n111_s;
                    stage6_col113[0] <= fa_s5_c112_n110_c;
                    stage6_col113[1] <= fa_s5_c112_n111_c;
                    stage6_col113[2] <= fa_s5_c113_n112_s;
                    stage6_col113[3] <= ha_s5_c113_n29_s;
                    stage6_col114[0] <= fa_s5_c113_n112_c;
                    stage6_col114[1] <= ha_s5_c113_n29_c;
                    stage6_col114[2] <= fa_s5_c114_n113_s;
                    stage6_col114[3] <= fa_s5_c114_n114_s;
                    stage6_col115[0] <= fa_s5_c114_n113_c;
                    stage6_col115[1] <= fa_s5_c114_n114_c;
                    stage6_col115[2] <= fa_s5_c115_n115_s;
                    stage6_col115[3] <= ha_s5_c115_n30_s;
                    stage6_col116[0] <= fa_s5_c115_n115_c;
                    stage6_col116[1] <= ha_s5_c115_n30_c;
                    stage6_col116[2] <= fa_s5_c116_n116_s;
                    stage6_col116[3] <= fa_s5_c116_n117_s;
                    stage6_col117[0] <= fa_s5_c116_n116_c;
                    stage6_col117[1] <= fa_s5_c116_n117_c;
                    stage6_col117[2] <= fa_s5_c117_n118_s;
                    stage6_col117[3] <= ha_s5_c117_n31_s;
                    stage6_col118[0] <= fa_s5_c117_n118_c;
                    stage6_col118[1] <= ha_s5_c117_n31_c;
                    stage6_col118[2] <= fa_s5_c118_n119_s;
                    stage6_col118[3] <= fa_s5_c118_n120_s;
                    stage6_col119[0] <= fa_s5_c118_n119_c;
                    stage6_col119[1] <= fa_s5_c118_n120_c;
                    stage6_col119[2] <= fa_s5_c119_n121_s;
                    stage6_col119[3] <= ha_s5_c119_n32_s;
                    stage6_col120[0] <= fa_s5_c119_n121_c;
                    stage6_col120[1] <= ha_s5_c119_n32_c;
                    stage6_col120[2] <= fa_s5_c120_n122_s;
                    stage6_col120[3] <= fa_s5_c120_n123_s;
                    stage6_col121[0] <= fa_s5_c120_n122_c;
                    stage6_col121[1] <= fa_s5_c120_n123_c;
                    stage6_col121[2] <= fa_s5_c121_n124_s;
                    stage6_col121[3] <= ha_s5_c121_n33_s;
                    stage6_col122[0] <= fa_s5_c121_n124_c;
                    stage6_col122[1] <= ha_s5_c121_n33_c;
                    stage6_col122[2] <= fa_s5_c122_n125_s;
                    stage6_col122[3] <= fa_s5_c122_n126_s;
                    stage6_col123[0] <= fa_s5_c122_n125_c;
                    stage6_col123[1] <= fa_s5_c122_n126_c;
                    stage6_col123[2] <= fa_s5_c123_n127_s;
                    stage6_col123[3] <= ha_s5_c123_n34_s;
                    stage6_col124[0] <= fa_s5_c123_n127_c;
                    stage6_col124[1] <= ha_s5_c123_n34_c;
                    stage6_col124[2] <= fa_s5_c124_n128_s;
                    stage6_col124[3] <= fa_s5_c124_n129_s;
                    stage6_col125[0] <= fa_s5_c124_n128_c;
                    stage6_col125[1] <= fa_s5_c124_n129_c;
                    stage6_col125[2] <= fa_s5_c125_n130_s;
                    stage6_col125[3] <= ha_s5_c125_n35_s;
                    stage6_col126[0] <= fa_s5_c125_n130_c;
                    stage6_col126[1] <= ha_s5_c125_n35_c;
                    stage6_col126[2] <= fa_s5_c126_n131_s;
                    stage6_col126[3] <= fa_s5_c126_n132_s;
                    stage6_col127[0] <= fa_s5_c126_n131_c;
                    stage6_col127[1] <= fa_s5_c126_n132_c;
                    stage6_col127[2] <= stage5_col127[0];
                    stage6_col127[3] <= stage5_col127[1];
                    stage6_col127[4] <= stage5_col127[2];
                    stage6_col127[5] <= stage5_col127[3];
                    stage6_col127[6] <= stage5_col127[4];
                    stage6_col127[7] <= stage5_col127[5];
                    stage6_col127[8] <= stage5_col127[6];
                    stage6_col127[9] <= stage5_col127[7];
                    stage6_col127[10] <= stage5_col127[8];
                    stage6_col127[11] <= stage5_col127[9];
                    stage6_col127[12] <= stage5_col127[10];
                    stage6_col127[13] <= stage5_col127[11];
                    stage6_col127[14] <= stage5_col127[12];
                    stage6_col127[15] <= stage5_col127[13];
                    stage6_col127[16] <= stage5_col127[14];
                    stage6_col127[17] <= stage5_col127[15];
                    stage6_col127[18] <= stage5_col127[16];
                    stage6_col127[19] <= stage5_col127[17];
                    stage6_col127[20] <= stage5_col127[18];
                    stage6_col127[21] <= stage5_col127[19];
                    stage6_col127[22] <= stage5_col127[20];
                    stage6_col127[23] <= stage5_col127[21];
                    stage6_col127[24] <= stage5_col127[22];
                    stage6_col127[25] <= stage5_col127[23];
                    stage6_col127[26] <= stage5_col127[24];
                    stage6_col127[27] <= stage5_col127[25];
                    stage6_col127[28] <= stage5_col127[26];
                    stage6_col127[29] <= stage5_col127[27];
                    stage6_col127[30] <= stage5_col127[27];
                    stage6_col127[31] <= stage5_col127[27];
                    stage6_col127[32] <= stage5_col127[27];
                    stage6_col127[33] <= stage5_col127[27];
                    stage6_col127[34] <= stage5_col127[27];
                    stage6_col127[35] <= stage5_col127[27];
                    stage6_col127[36] <= stage5_col127[27];
                    stage6_col127[37] <= stage5_col127[27];
                    stage6_col127[38] <= stage5_col127[27];
                    stage6_col127[39] <= stage5_col127[27];
                    stage6_col127[40] <= stage5_col127[27];
                    stage6_col127[41] <= stage5_col127[27];
                    stage6_col127[42] <= stage5_col127[27];
                    stage6_col127[43] <= stage5_col127[27];
                    stage6_col127[44] <= stage5_col127[27];
                    stage6_col127[45] <= stage5_col127[27];
                    stage6_col127[46] <= stage5_col127[27];
                    stage6_col127[47] <= stage5_col127[27];
                    stage6_col127[48] <= stage5_col127[27];
                    stage6_col127[49] <= stage5_col127[27];
                    stage6_col127[50] <= stage5_col127[27];
                    stage6_col127[51] <= stage5_col127[27];
                    stage6_col127[52] <= stage5_col127[27];
                    stage6_col127[53] <= stage5_col127[27];
                    stage6_col127[54] <= stage5_col127[27];
                    stage6_col127[55] <= stage5_col127[27];
                    stage6_col127[56] <= stage5_col127[27];
                    stage6_col127[57] <= stage5_col127[27];
                    stage6_col127[58] <= stage5_col127[27];
                    stage6_col127[59] <= stage5_col127[27];
                    stage6_col127[60] <= stage5_col127[27];
                end
            end
        end else begin : gen_stage6_no_pipe
            // Combinational assignment
            always_comb begin
                stage6_col0[0] = stage5_col0[0];
                stage6_col1[0] = stage5_col1[0];
                stage6_col2[0] = stage5_col2[0];
                stage6_col3[0] = stage5_col3[0];
                stage6_col4[0] = stage5_col4[0];
                stage6_col5[0] = ha_s5_c5_n0_s;
                stage6_col6[0] = ha_s5_c5_n0_c;
                stage6_col6[1] = stage5_col6[0];
                stage6_col7[0] = fa_s5_c7_n0_s;
                stage6_col8[0] = fa_s5_c7_n0_c;
                stage6_col8[1] = stage5_col8[0];
                stage6_col8[2] = stage5_col8[1];
                stage6_col9[0] = stage5_col9[0];
                stage6_col9[1] = stage5_col9[1];
                stage6_col10[0] = stage5_col10[0];
                stage6_col10[1] = stage5_col10[1];
                stage6_col11[0] = stage5_col11[0];
                stage6_col11[1] = stage5_col11[1];
                stage6_col12[0] = stage5_col12[0];
                stage6_col12[1] = stage5_col12[1];
                stage6_col13[0] = stage5_col13[0];
                stage6_col13[1] = stage5_col13[1];
                stage6_col14[0] = stage5_col14[0];
                stage6_col14[1] = stage5_col14[1];
                stage6_col15[0] = stage5_col15[0];
                stage6_col15[1] = stage5_col15[1];
                stage6_col16[0] = stage5_col16[0];
                stage6_col16[1] = stage5_col16[1];
                stage6_col17[0] = stage5_col17[0];
                stage6_col17[1] = stage5_col17[1];
                stage6_col18[0] = stage5_col18[0];
                stage6_col18[1] = stage5_col18[1];
                stage6_col19[0] = stage5_col19[0];
                stage6_col19[1] = stage5_col19[1];
                stage6_col20[0] = stage5_col20[0];
                stage6_col20[1] = stage5_col20[1];
                stage6_col21[0] = stage5_col21[0];
                stage6_col21[1] = stage5_col21[1];
                stage6_col22[0] = stage5_col22[0];
                stage6_col22[1] = stage5_col22[1];
                stage6_col23[0] = stage5_col23[0];
                stage6_col23[1] = stage5_col23[1];
                stage6_col24[0] = stage5_col24[0];
                stage6_col24[1] = stage5_col24[1];
                stage6_col25[0] = stage5_col25[0];
                stage6_col25[1] = stage5_col25[1];
                stage6_col26[0] = stage5_col26[0];
                stage6_col26[1] = stage5_col26[1];
                stage6_col27[0] = stage5_col27[0];
                stage6_col27[1] = stage5_col27[1];
                stage6_col28[0] = fa_s5_c28_n1_s;
                stage6_col28[1] = stage5_col28[3];
                stage6_col29[0] = fa_s5_c28_n1_c;
                stage6_col29[1] = fa_s5_c29_n2_s;
                stage6_col30[0] = fa_s5_c29_n2_c;
                stage6_col30[1] = fa_s5_c30_n3_s;
                stage6_col31[0] = fa_s5_c30_n3_c;
                stage6_col31[1] = fa_s5_c31_n4_s;
                stage6_col32[0] = fa_s5_c31_n4_c;
                stage6_col32[1] = fa_s5_c32_n5_s;
                stage6_col33[0] = fa_s5_c32_n5_c;
                stage6_col33[1] = fa_s5_c33_n6_s;
                stage6_col34[0] = fa_s5_c33_n6_c;
                stage6_col34[1] = fa_s5_c34_n7_s;
                stage6_col35[0] = fa_s5_c34_n7_c;
                stage6_col35[1] = fa_s5_c35_n8_s;
                stage6_col36[0] = fa_s5_c35_n8_c;
                stage6_col36[1] = fa_s5_c36_n9_s;
                stage6_col37[0] = fa_s5_c36_n9_c;
                stage6_col37[1] = fa_s5_c37_n10_s;
                stage6_col38[0] = fa_s5_c37_n10_c;
                stage6_col38[1] = fa_s5_c38_n11_s;
                stage6_col39[0] = fa_s5_c38_n11_c;
                stage6_col39[1] = fa_s5_c39_n12_s;
                stage6_col40[0] = fa_s5_c39_n12_c;
                stage6_col40[1] = fa_s5_c40_n13_s;
                stage6_col41[0] = fa_s5_c40_n13_c;
                stage6_col41[1] = fa_s5_c41_n14_s;
                stage6_col41[2] = stage5_col41[3];
                stage6_col41[3] = stage5_col41[4];
                stage6_col42[0] = fa_s5_c41_n14_c;
                stage6_col42[1] = fa_s5_c42_n15_s;
                stage6_col42[2] = stage5_col42[3];
                stage6_col43[0] = fa_s5_c42_n15_c;
                stage6_col43[1] = fa_s5_c43_n16_s;
                stage6_col43[2] = stage5_col43[3];
                stage6_col44[0] = fa_s5_c43_n16_c;
                stage6_col44[1] = fa_s5_c44_n17_s;
                stage6_col44[2] = stage5_col44[3];
                stage6_col45[0] = fa_s5_c44_n17_c;
                stage6_col45[1] = fa_s5_c45_n18_s;
                stage6_col45[2] = stage5_col45[3];
                stage6_col46[0] = fa_s5_c45_n18_c;
                stage6_col46[1] = fa_s5_c46_n19_s;
                stage6_col46[2] = stage5_col46[3];
                stage6_col47[0] = fa_s5_c46_n19_c;
                stage6_col47[1] = fa_s5_c47_n20_s;
                stage6_col47[2] = stage5_col47[3];
                stage6_col48[0] = fa_s5_c47_n20_c;
                stage6_col48[1] = fa_s5_c48_n21_s;
                stage6_col48[2] = stage5_col48[3];
                stage6_col49[0] = fa_s5_c48_n21_c;
                stage6_col49[1] = fa_s5_c49_n22_s;
                stage6_col49[2] = stage5_col49[3];
                stage6_col50[0] = fa_s5_c49_n22_c;
                stage6_col50[1] = fa_s5_c50_n23_s;
                stage6_col50[2] = stage5_col50[3];
                stage6_col51[0] = fa_s5_c50_n23_c;
                stage6_col51[1] = fa_s5_c51_n24_s;
                stage6_col51[2] = stage5_col51[3];
                stage6_col52[0] = fa_s5_c51_n24_c;
                stage6_col52[1] = fa_s5_c52_n25_s;
                stage6_col52[2] = stage5_col52[3];
                stage6_col53[0] = fa_s5_c52_n25_c;
                stage6_col53[1] = fa_s5_c53_n26_s;
                stage6_col53[2] = stage5_col53[3];
                stage6_col54[0] = fa_s5_c53_n26_c;
                stage6_col54[1] = fa_s5_c54_n27_s;
                stage6_col54[2] = stage5_col54[3];
                stage6_col55[0] = fa_s5_c54_n27_c;
                stage6_col55[1] = fa_s5_c55_n28_s;
                stage6_col55[2] = stage5_col55[3];
                stage6_col56[0] = fa_s5_c55_n28_c;
                stage6_col56[1] = fa_s5_c56_n29_s;
                stage6_col56[2] = stage5_col56[3];
                stage6_col57[0] = fa_s5_c56_n29_c;
                stage6_col57[1] = fa_s5_c57_n30_s;
                stage6_col57[2] = stage5_col57[3];
                stage6_col58[0] = fa_s5_c57_n30_c;
                stage6_col58[1] = fa_s5_c58_n31_s;
                stage6_col58[2] = stage5_col58[3];
                stage6_col59[0] = fa_s5_c58_n31_c;
                stage6_col59[1] = fa_s5_c59_n32_s;
                stage6_col59[2] = fa_s5_c59_n33_s;
                stage6_col60[0] = fa_s5_c59_n32_c;
                stage6_col60[1] = fa_s5_c59_n33_c;
                stage6_col60[2] = fa_s5_c60_n34_s;
                stage6_col60[3] = ha_s5_c60_n1_s;
                stage6_col61[0] = fa_s5_c60_n34_c;
                stage6_col61[1] = ha_s5_c60_n1_c;
                stage6_col61[2] = fa_s5_c61_n35_s;
                stage6_col61[3] = ha_s5_c61_n2_s;
                stage6_col62[0] = fa_s5_c61_n35_c;
                stage6_col62[1] = ha_s5_c61_n2_c;
                stage6_col62[2] = fa_s5_c62_n36_s;
                stage6_col62[3] = ha_s5_c62_n3_s;
                stage6_col63[0] = fa_s5_c62_n36_c;
                stage6_col63[1] = ha_s5_c62_n3_c;
                stage6_col63[2] = fa_s5_c63_n37_s;
                stage6_col63[3] = ha_s5_c63_n4_s;
                stage6_col64[0] = fa_s5_c63_n37_c;
                stage6_col64[1] = ha_s5_c63_n4_c;
                stage6_col64[2] = fa_s5_c64_n38_s;
                stage6_col64[3] = fa_s5_c64_n39_s;
                stage6_col65[0] = fa_s5_c64_n38_c;
                stage6_col65[1] = fa_s5_c64_n39_c;
                stage6_col65[2] = fa_s5_c65_n40_s;
                stage6_col65[3] = ha_s5_c65_n5_s;
                stage6_col66[0] = fa_s5_c65_n40_c;
                stage6_col66[1] = ha_s5_c65_n5_c;
                stage6_col66[2] = fa_s5_c66_n41_s;
                stage6_col66[3] = fa_s5_c66_n42_s;
                stage6_col67[0] = fa_s5_c66_n41_c;
                stage6_col67[1] = fa_s5_c66_n42_c;
                stage6_col67[2] = fa_s5_c67_n43_s;
                stage6_col67[3] = ha_s5_c67_n6_s;
                stage6_col68[0] = fa_s5_c67_n43_c;
                stage6_col68[1] = ha_s5_c67_n6_c;
                stage6_col68[2] = fa_s5_c68_n44_s;
                stage6_col68[3] = fa_s5_c68_n45_s;
                stage6_col69[0] = fa_s5_c68_n44_c;
                stage6_col69[1] = fa_s5_c68_n45_c;
                stage6_col69[2] = fa_s5_c69_n46_s;
                stage6_col69[3] = ha_s5_c69_n7_s;
                stage6_col70[0] = fa_s5_c69_n46_c;
                stage6_col70[1] = ha_s5_c69_n7_c;
                stage6_col70[2] = fa_s5_c70_n47_s;
                stage6_col70[3] = fa_s5_c70_n48_s;
                stage6_col71[0] = fa_s5_c70_n47_c;
                stage6_col71[1] = fa_s5_c70_n48_c;
                stage6_col71[2] = fa_s5_c71_n49_s;
                stage6_col71[3] = ha_s5_c71_n8_s;
                stage6_col72[0] = fa_s5_c71_n49_c;
                stage6_col72[1] = ha_s5_c71_n8_c;
                stage6_col72[2] = fa_s5_c72_n50_s;
                stage6_col72[3] = fa_s5_c72_n51_s;
                stage6_col73[0] = fa_s5_c72_n50_c;
                stage6_col73[1] = fa_s5_c72_n51_c;
                stage6_col73[2] = fa_s5_c73_n52_s;
                stage6_col73[3] = ha_s5_c73_n9_s;
                stage6_col74[0] = fa_s5_c73_n52_c;
                stage6_col74[1] = ha_s5_c73_n9_c;
                stage6_col74[2] = fa_s5_c74_n53_s;
                stage6_col74[3] = fa_s5_c74_n54_s;
                stage6_col75[0] = fa_s5_c74_n53_c;
                stage6_col75[1] = fa_s5_c74_n54_c;
                stage6_col75[2] = fa_s5_c75_n55_s;
                stage6_col75[3] = ha_s5_c75_n10_s;
                stage6_col76[0] = fa_s5_c75_n55_c;
                stage6_col76[1] = ha_s5_c75_n10_c;
                stage6_col76[2] = fa_s5_c76_n56_s;
                stage6_col76[3] = fa_s5_c76_n57_s;
                stage6_col77[0] = fa_s5_c76_n56_c;
                stage6_col77[1] = fa_s5_c76_n57_c;
                stage6_col77[2] = fa_s5_c77_n58_s;
                stage6_col77[3] = ha_s5_c77_n11_s;
                stage6_col78[0] = fa_s5_c77_n58_c;
                stage6_col78[1] = ha_s5_c77_n11_c;
                stage6_col78[2] = fa_s5_c78_n59_s;
                stage6_col78[3] = fa_s5_c78_n60_s;
                stage6_col79[0] = fa_s5_c78_n59_c;
                stage6_col79[1] = fa_s5_c78_n60_c;
                stage6_col79[2] = fa_s5_c79_n61_s;
                stage6_col79[3] = ha_s5_c79_n12_s;
                stage6_col80[0] = fa_s5_c79_n61_c;
                stage6_col80[1] = ha_s5_c79_n12_c;
                stage6_col80[2] = fa_s5_c80_n62_s;
                stage6_col80[3] = fa_s5_c80_n63_s;
                stage6_col81[0] = fa_s5_c80_n62_c;
                stage6_col81[1] = fa_s5_c80_n63_c;
                stage6_col81[2] = fa_s5_c81_n64_s;
                stage6_col81[3] = ha_s5_c81_n13_s;
                stage6_col82[0] = fa_s5_c81_n64_c;
                stage6_col82[1] = ha_s5_c81_n13_c;
                stage6_col82[2] = fa_s5_c82_n65_s;
                stage6_col82[3] = fa_s5_c82_n66_s;
                stage6_col83[0] = fa_s5_c82_n65_c;
                stage6_col83[1] = fa_s5_c82_n66_c;
                stage6_col83[2] = fa_s5_c83_n67_s;
                stage6_col83[3] = ha_s5_c83_n14_s;
                stage6_col84[0] = fa_s5_c83_n67_c;
                stage6_col84[1] = ha_s5_c83_n14_c;
                stage6_col84[2] = fa_s5_c84_n68_s;
                stage6_col84[3] = fa_s5_c84_n69_s;
                stage6_col85[0] = fa_s5_c84_n68_c;
                stage6_col85[1] = fa_s5_c84_n69_c;
                stage6_col85[2] = fa_s5_c85_n70_s;
                stage6_col85[3] = ha_s5_c85_n15_s;
                stage6_col86[0] = fa_s5_c85_n70_c;
                stage6_col86[1] = ha_s5_c85_n15_c;
                stage6_col86[2] = fa_s5_c86_n71_s;
                stage6_col86[3] = fa_s5_c86_n72_s;
                stage6_col87[0] = fa_s5_c86_n71_c;
                stage6_col87[1] = fa_s5_c86_n72_c;
                stage6_col87[2] = fa_s5_c87_n73_s;
                stage6_col87[3] = ha_s5_c87_n16_s;
                stage6_col88[0] = fa_s5_c87_n73_c;
                stage6_col88[1] = ha_s5_c87_n16_c;
                stage6_col88[2] = fa_s5_c88_n74_s;
                stage6_col88[3] = fa_s5_c88_n75_s;
                stage6_col89[0] = fa_s5_c88_n74_c;
                stage6_col89[1] = fa_s5_c88_n75_c;
                stage6_col89[2] = fa_s5_c89_n76_s;
                stage6_col89[3] = ha_s5_c89_n17_s;
                stage6_col90[0] = fa_s5_c89_n76_c;
                stage6_col90[1] = ha_s5_c89_n17_c;
                stage6_col90[2] = fa_s5_c90_n77_s;
                stage6_col90[3] = fa_s5_c90_n78_s;
                stage6_col91[0] = fa_s5_c90_n77_c;
                stage6_col91[1] = fa_s5_c90_n78_c;
                stage6_col91[2] = fa_s5_c91_n79_s;
                stage6_col91[3] = ha_s5_c91_n18_s;
                stage6_col92[0] = fa_s5_c91_n79_c;
                stage6_col92[1] = ha_s5_c91_n18_c;
                stage6_col92[2] = fa_s5_c92_n80_s;
                stage6_col92[3] = fa_s5_c92_n81_s;
                stage6_col93[0] = fa_s5_c92_n80_c;
                stage6_col93[1] = fa_s5_c92_n81_c;
                stage6_col93[2] = fa_s5_c93_n82_s;
                stage6_col93[3] = ha_s5_c93_n19_s;
                stage6_col94[0] = fa_s5_c93_n82_c;
                stage6_col94[1] = ha_s5_c93_n19_c;
                stage6_col94[2] = fa_s5_c94_n83_s;
                stage6_col94[3] = fa_s5_c94_n84_s;
                stage6_col95[0] = fa_s5_c94_n83_c;
                stage6_col95[1] = fa_s5_c94_n84_c;
                stage6_col95[2] = fa_s5_c95_n85_s;
                stage6_col95[3] = ha_s5_c95_n20_s;
                stage6_col96[0] = fa_s5_c95_n85_c;
                stage6_col96[1] = ha_s5_c95_n20_c;
                stage6_col96[2] = fa_s5_c96_n86_s;
                stage6_col96[3] = fa_s5_c96_n87_s;
                stage6_col97[0] = fa_s5_c96_n86_c;
                stage6_col97[1] = fa_s5_c96_n87_c;
                stage6_col97[2] = fa_s5_c97_n88_s;
                stage6_col97[3] = ha_s5_c97_n21_s;
                stage6_col98[0] = fa_s5_c97_n88_c;
                stage6_col98[1] = ha_s5_c97_n21_c;
                stage6_col98[2] = fa_s5_c98_n89_s;
                stage6_col98[3] = fa_s5_c98_n90_s;
                stage6_col99[0] = fa_s5_c98_n89_c;
                stage6_col99[1] = fa_s5_c98_n90_c;
                stage6_col99[2] = fa_s5_c99_n91_s;
                stage6_col99[3] = ha_s5_c99_n22_s;
                stage6_col100[0] = fa_s5_c99_n91_c;
                stage6_col100[1] = ha_s5_c99_n22_c;
                stage6_col100[2] = fa_s5_c100_n92_s;
                stage6_col100[3] = fa_s5_c100_n93_s;
                stage6_col101[0] = fa_s5_c100_n92_c;
                stage6_col101[1] = fa_s5_c100_n93_c;
                stage6_col101[2] = fa_s5_c101_n94_s;
                stage6_col101[3] = ha_s5_c101_n23_s;
                stage6_col102[0] = fa_s5_c101_n94_c;
                stage6_col102[1] = ha_s5_c101_n23_c;
                stage6_col102[2] = fa_s5_c102_n95_s;
                stage6_col102[3] = fa_s5_c102_n96_s;
                stage6_col103[0] = fa_s5_c102_n95_c;
                stage6_col103[1] = fa_s5_c102_n96_c;
                stage6_col103[2] = fa_s5_c103_n97_s;
                stage6_col103[3] = ha_s5_c103_n24_s;
                stage6_col104[0] = fa_s5_c103_n97_c;
                stage6_col104[1] = ha_s5_c103_n24_c;
                stage6_col104[2] = fa_s5_c104_n98_s;
                stage6_col104[3] = fa_s5_c104_n99_s;
                stage6_col105[0] = fa_s5_c104_n98_c;
                stage6_col105[1] = fa_s5_c104_n99_c;
                stage6_col105[2] = fa_s5_c105_n100_s;
                stage6_col105[3] = ha_s5_c105_n25_s;
                stage6_col106[0] = fa_s5_c105_n100_c;
                stage6_col106[1] = ha_s5_c105_n25_c;
                stage6_col106[2] = fa_s5_c106_n101_s;
                stage6_col106[3] = fa_s5_c106_n102_s;
                stage6_col107[0] = fa_s5_c106_n101_c;
                stage6_col107[1] = fa_s5_c106_n102_c;
                stage6_col107[2] = fa_s5_c107_n103_s;
                stage6_col107[3] = ha_s5_c107_n26_s;
                stage6_col108[0] = fa_s5_c107_n103_c;
                stage6_col108[1] = ha_s5_c107_n26_c;
                stage6_col108[2] = fa_s5_c108_n104_s;
                stage6_col108[3] = fa_s5_c108_n105_s;
                stage6_col109[0] = fa_s5_c108_n104_c;
                stage6_col109[1] = fa_s5_c108_n105_c;
                stage6_col109[2] = fa_s5_c109_n106_s;
                stage6_col109[3] = ha_s5_c109_n27_s;
                stage6_col110[0] = fa_s5_c109_n106_c;
                stage6_col110[1] = ha_s5_c109_n27_c;
                stage6_col110[2] = fa_s5_c110_n107_s;
                stage6_col110[3] = fa_s5_c110_n108_s;
                stage6_col111[0] = fa_s5_c110_n107_c;
                stage6_col111[1] = fa_s5_c110_n108_c;
                stage6_col111[2] = fa_s5_c111_n109_s;
                stage6_col111[3] = ha_s5_c111_n28_s;
                stage6_col112[0] = fa_s5_c111_n109_c;
                stage6_col112[1] = ha_s5_c111_n28_c;
                stage6_col112[2] = fa_s5_c112_n110_s;
                stage6_col112[3] = fa_s5_c112_n111_s;
                stage6_col113[0] = fa_s5_c112_n110_c;
                stage6_col113[1] = fa_s5_c112_n111_c;
                stage6_col113[2] = fa_s5_c113_n112_s;
                stage6_col113[3] = ha_s5_c113_n29_s;
                stage6_col114[0] = fa_s5_c113_n112_c;
                stage6_col114[1] = ha_s5_c113_n29_c;
                stage6_col114[2] = fa_s5_c114_n113_s;
                stage6_col114[3] = fa_s5_c114_n114_s;
                stage6_col115[0] = fa_s5_c114_n113_c;
                stage6_col115[1] = fa_s5_c114_n114_c;
                stage6_col115[2] = fa_s5_c115_n115_s;
                stage6_col115[3] = ha_s5_c115_n30_s;
                stage6_col116[0] = fa_s5_c115_n115_c;
                stage6_col116[1] = ha_s5_c115_n30_c;
                stage6_col116[2] = fa_s5_c116_n116_s;
                stage6_col116[3] = fa_s5_c116_n117_s;
                stage6_col117[0] = fa_s5_c116_n116_c;
                stage6_col117[1] = fa_s5_c116_n117_c;
                stage6_col117[2] = fa_s5_c117_n118_s;
                stage6_col117[3] = ha_s5_c117_n31_s;
                stage6_col118[0] = fa_s5_c117_n118_c;
                stage6_col118[1] = ha_s5_c117_n31_c;
                stage6_col118[2] = fa_s5_c118_n119_s;
                stage6_col118[3] = fa_s5_c118_n120_s;
                stage6_col119[0] = fa_s5_c118_n119_c;
                stage6_col119[1] = fa_s5_c118_n120_c;
                stage6_col119[2] = fa_s5_c119_n121_s;
                stage6_col119[3] = ha_s5_c119_n32_s;
                stage6_col120[0] = fa_s5_c119_n121_c;
                stage6_col120[1] = ha_s5_c119_n32_c;
                stage6_col120[2] = fa_s5_c120_n122_s;
                stage6_col120[3] = fa_s5_c120_n123_s;
                stage6_col121[0] = fa_s5_c120_n122_c;
                stage6_col121[1] = fa_s5_c120_n123_c;
                stage6_col121[2] = fa_s5_c121_n124_s;
                stage6_col121[3] = ha_s5_c121_n33_s;
                stage6_col122[0] = fa_s5_c121_n124_c;
                stage6_col122[1] = ha_s5_c121_n33_c;
                stage6_col122[2] = fa_s5_c122_n125_s;
                stage6_col122[3] = fa_s5_c122_n126_s;
                stage6_col123[0] = fa_s5_c122_n125_c;
                stage6_col123[1] = fa_s5_c122_n126_c;
                stage6_col123[2] = fa_s5_c123_n127_s;
                stage6_col123[3] = ha_s5_c123_n34_s;
                stage6_col124[0] = fa_s5_c123_n127_c;
                stage6_col124[1] = ha_s5_c123_n34_c;
                stage6_col124[2] = fa_s5_c124_n128_s;
                stage6_col124[3] = fa_s5_c124_n129_s;
                stage6_col125[0] = fa_s5_c124_n128_c;
                stage6_col125[1] = fa_s5_c124_n129_c;
                stage6_col125[2] = fa_s5_c125_n130_s;
                stage6_col125[3] = ha_s5_c125_n35_s;
                stage6_col126[0] = fa_s5_c125_n130_c;
                stage6_col126[1] = ha_s5_c125_n35_c;
                stage6_col126[2] = fa_s5_c126_n131_s;
                stage6_col126[3] = fa_s5_c126_n132_s;
                stage6_col127[0] = fa_s5_c126_n131_c;
                stage6_col127[1] = fa_s5_c126_n132_c;
                stage6_col127[2] = stage5_col127[0];
                stage6_col127[3] = stage5_col127[1];
                stage6_col127[4] = stage5_col127[2];
                stage6_col127[5] = stage5_col127[3];
                stage6_col127[6] = stage5_col127[4];
                stage6_col127[7] = stage5_col127[5];
                stage6_col127[8] = stage5_col127[6];
                stage6_col127[9] = stage5_col127[7];
                stage6_col127[10] = stage5_col127[8];
                stage6_col127[11] = stage5_col127[9];
                stage6_col127[12] = stage5_col127[10];
                stage6_col127[13] = stage5_col127[11];
                stage6_col127[14] = stage5_col127[12];
                stage6_col127[15] = stage5_col127[13];
                stage6_col127[16] = stage5_col127[14];
                stage6_col127[17] = stage5_col127[15];
                stage6_col127[18] = stage5_col127[16];
                stage6_col127[19] = stage5_col127[17];
                stage6_col127[20] = stage5_col127[18];
                stage6_col127[21] = stage5_col127[19];
                stage6_col127[22] = stage5_col127[20];
                stage6_col127[23] = stage5_col127[21];
                stage6_col127[24] = stage5_col127[22];
                stage6_col127[25] = stage5_col127[23];
                stage6_col127[26] = stage5_col127[24];
                stage6_col127[27] = stage5_col127[25];
                stage6_col127[28] = stage5_col127[26];
                stage6_col127[29] = stage5_col127[27];
                stage6_col127[30] = stage5_col127[27];
                stage6_col127[31] = stage5_col127[27];
                stage6_col127[32] = stage5_col127[27];
                stage6_col127[33] = stage5_col127[27];
                stage6_col127[34] = stage5_col127[27];
                stage6_col127[35] = stage5_col127[27];
                stage6_col127[36] = stage5_col127[27];
                stage6_col127[37] = stage5_col127[27];
                stage6_col127[38] = stage5_col127[27];
                stage6_col127[39] = stage5_col127[27];
                stage6_col127[40] = stage5_col127[27];
                stage6_col127[41] = stage5_col127[27];
                stage6_col127[42] = stage5_col127[27];
                stage6_col127[43] = stage5_col127[27];
                stage6_col127[44] = stage5_col127[27];
                stage6_col127[45] = stage5_col127[27];
                stage6_col127[46] = stage5_col127[27];
                stage6_col127[47] = stage5_col127[27];
                stage6_col127[48] = stage5_col127[27];
                stage6_col127[49] = stage5_col127[27];
                stage6_col127[50] = stage5_col127[27];
                stage6_col127[51] = stage5_col127[27];
                stage6_col127[52] = stage5_col127[27];
                stage6_col127[53] = stage5_col127[27];
                stage6_col127[54] = stage5_col127[27];
                stage6_col127[55] = stage5_col127[27];
                stage6_col127[56] = stage5_col127[27];
                stage6_col127[57] = stage5_col127[27];
                stage6_col127[58] = stage5_col127[27];
                stage6_col127[59] = stage5_col127[27];
                stage6_col127[60] = stage5_col127[27];
            end
        end
    endgenerate

    // Stage 7: Reduction
    fa fa_s6_c8_n0 (
        .a(stage6_col8[0]),
        .b(stage6_col8[1]),
        .c_in(stage6_col8[2]),
        .s(fa_s6_c8_n0_s),
        .c_out(fa_s6_c8_n0_c)
    );

    fa fa_s6_c41_n1 (
        .a(stage6_col41[0]),
        .b(stage6_col41[1]),
        .c_in(stage6_col41[2]),
        .s(fa_s6_c41_n1_s),
        .c_out(fa_s6_c41_n1_c)
    );

    fa fa_s6_c42_n2 (
        .a(stage6_col42[0]),
        .b(stage6_col42[1]),
        .c_in(stage6_col42[2]),
        .s(fa_s6_c42_n2_s),
        .c_out(fa_s6_c42_n2_c)
    );

    fa fa_s6_c43_n3 (
        .a(stage6_col43[0]),
        .b(stage6_col43[1]),
        .c_in(stage6_col43[2]),
        .s(fa_s6_c43_n3_s),
        .c_out(fa_s6_c43_n3_c)
    );

    fa fa_s6_c44_n4 (
        .a(stage6_col44[0]),
        .b(stage6_col44[1]),
        .c_in(stage6_col44[2]),
        .s(fa_s6_c44_n4_s),
        .c_out(fa_s6_c44_n4_c)
    );

    fa fa_s6_c45_n5 (
        .a(stage6_col45[0]),
        .b(stage6_col45[1]),
        .c_in(stage6_col45[2]),
        .s(fa_s6_c45_n5_s),
        .c_out(fa_s6_c45_n5_c)
    );

    fa fa_s6_c46_n6 (
        .a(stage6_col46[0]),
        .b(stage6_col46[1]),
        .c_in(stage6_col46[2]),
        .s(fa_s6_c46_n6_s),
        .c_out(fa_s6_c46_n6_c)
    );

    fa fa_s6_c47_n7 (
        .a(stage6_col47[0]),
        .b(stage6_col47[1]),
        .c_in(stage6_col47[2]),
        .s(fa_s6_c47_n7_s),
        .c_out(fa_s6_c47_n7_c)
    );

    fa fa_s6_c48_n8 (
        .a(stage6_col48[0]),
        .b(stage6_col48[1]),
        .c_in(stage6_col48[2]),
        .s(fa_s6_c48_n8_s),
        .c_out(fa_s6_c48_n8_c)
    );

    fa fa_s6_c49_n9 (
        .a(stage6_col49[0]),
        .b(stage6_col49[1]),
        .c_in(stage6_col49[2]),
        .s(fa_s6_c49_n9_s),
        .c_out(fa_s6_c49_n9_c)
    );

    fa fa_s6_c50_n10 (
        .a(stage6_col50[0]),
        .b(stage6_col50[1]),
        .c_in(stage6_col50[2]),
        .s(fa_s6_c50_n10_s),
        .c_out(fa_s6_c50_n10_c)
    );

    fa fa_s6_c51_n11 (
        .a(stage6_col51[0]),
        .b(stage6_col51[1]),
        .c_in(stage6_col51[2]),
        .s(fa_s6_c51_n11_s),
        .c_out(fa_s6_c51_n11_c)
    );

    fa fa_s6_c52_n12 (
        .a(stage6_col52[0]),
        .b(stage6_col52[1]),
        .c_in(stage6_col52[2]),
        .s(fa_s6_c52_n12_s),
        .c_out(fa_s6_c52_n12_c)
    );

    fa fa_s6_c53_n13 (
        .a(stage6_col53[0]),
        .b(stage6_col53[1]),
        .c_in(stage6_col53[2]),
        .s(fa_s6_c53_n13_s),
        .c_out(fa_s6_c53_n13_c)
    );

    fa fa_s6_c54_n14 (
        .a(stage6_col54[0]),
        .b(stage6_col54[1]),
        .c_in(stage6_col54[2]),
        .s(fa_s6_c54_n14_s),
        .c_out(fa_s6_c54_n14_c)
    );

    fa fa_s6_c55_n15 (
        .a(stage6_col55[0]),
        .b(stage6_col55[1]),
        .c_in(stage6_col55[2]),
        .s(fa_s6_c55_n15_s),
        .c_out(fa_s6_c55_n15_c)
    );

    fa fa_s6_c56_n16 (
        .a(stage6_col56[0]),
        .b(stage6_col56[1]),
        .c_in(stage6_col56[2]),
        .s(fa_s6_c56_n16_s),
        .c_out(fa_s6_c56_n16_c)
    );

    fa fa_s6_c57_n17 (
        .a(stage6_col57[0]),
        .b(stage6_col57[1]),
        .c_in(stage6_col57[2]),
        .s(fa_s6_c57_n17_s),
        .c_out(fa_s6_c57_n17_c)
    );

    fa fa_s6_c58_n18 (
        .a(stage6_col58[0]),
        .b(stage6_col58[1]),
        .c_in(stage6_col58[2]),
        .s(fa_s6_c58_n18_s),
        .c_out(fa_s6_c58_n18_c)
    );

    fa fa_s6_c59_n19 (
        .a(stage6_col59[0]),
        .b(stage6_col59[1]),
        .c_in(stage6_col59[2]),
        .s(fa_s6_c59_n19_s),
        .c_out(fa_s6_c59_n19_c)
    );

    fa fa_s6_c60_n20 (
        .a(stage6_col60[0]),
        .b(stage6_col60[1]),
        .c_in(stage6_col60[2]),
        .s(fa_s6_c60_n20_s),
        .c_out(fa_s6_c60_n20_c)
    );

    fa fa_s6_c61_n21 (
        .a(stage6_col61[0]),
        .b(stage6_col61[1]),
        .c_in(stage6_col61[2]),
        .s(fa_s6_c61_n21_s),
        .c_out(fa_s6_c61_n21_c)
    );

    fa fa_s6_c62_n22 (
        .a(stage6_col62[0]),
        .b(stage6_col62[1]),
        .c_in(stage6_col62[2]),
        .s(fa_s6_c62_n22_s),
        .c_out(fa_s6_c62_n22_c)
    );

    fa fa_s6_c63_n23 (
        .a(stage6_col63[0]),
        .b(stage6_col63[1]),
        .c_in(stage6_col63[2]),
        .s(fa_s6_c63_n23_s),
        .c_out(fa_s6_c63_n23_c)
    );

    fa fa_s6_c64_n24 (
        .a(stage6_col64[0]),
        .b(stage6_col64[1]),
        .c_in(stage6_col64[2]),
        .s(fa_s6_c64_n24_s),
        .c_out(fa_s6_c64_n24_c)
    );

    fa fa_s6_c65_n25 (
        .a(stage6_col65[0]),
        .b(stage6_col65[1]),
        .c_in(stage6_col65[2]),
        .s(fa_s6_c65_n25_s),
        .c_out(fa_s6_c65_n25_c)
    );

    fa fa_s6_c66_n26 (
        .a(stage6_col66[0]),
        .b(stage6_col66[1]),
        .c_in(stage6_col66[2]),
        .s(fa_s6_c66_n26_s),
        .c_out(fa_s6_c66_n26_c)
    );

    fa fa_s6_c67_n27 (
        .a(stage6_col67[0]),
        .b(stage6_col67[1]),
        .c_in(stage6_col67[2]),
        .s(fa_s6_c67_n27_s),
        .c_out(fa_s6_c67_n27_c)
    );

    fa fa_s6_c68_n28 (
        .a(stage6_col68[0]),
        .b(stage6_col68[1]),
        .c_in(stage6_col68[2]),
        .s(fa_s6_c68_n28_s),
        .c_out(fa_s6_c68_n28_c)
    );

    fa fa_s6_c69_n29 (
        .a(stage6_col69[0]),
        .b(stage6_col69[1]),
        .c_in(stage6_col69[2]),
        .s(fa_s6_c69_n29_s),
        .c_out(fa_s6_c69_n29_c)
    );

    fa fa_s6_c70_n30 (
        .a(stage6_col70[0]),
        .b(stage6_col70[1]),
        .c_in(stage6_col70[2]),
        .s(fa_s6_c70_n30_s),
        .c_out(fa_s6_c70_n30_c)
    );

    fa fa_s6_c71_n31 (
        .a(stage6_col71[0]),
        .b(stage6_col71[1]),
        .c_in(stage6_col71[2]),
        .s(fa_s6_c71_n31_s),
        .c_out(fa_s6_c71_n31_c)
    );

    fa fa_s6_c72_n32 (
        .a(stage6_col72[0]),
        .b(stage6_col72[1]),
        .c_in(stage6_col72[2]),
        .s(fa_s6_c72_n32_s),
        .c_out(fa_s6_c72_n32_c)
    );

    fa fa_s6_c73_n33 (
        .a(stage6_col73[0]),
        .b(stage6_col73[1]),
        .c_in(stage6_col73[2]),
        .s(fa_s6_c73_n33_s),
        .c_out(fa_s6_c73_n33_c)
    );

    fa fa_s6_c74_n34 (
        .a(stage6_col74[0]),
        .b(stage6_col74[1]),
        .c_in(stage6_col74[2]),
        .s(fa_s6_c74_n34_s),
        .c_out(fa_s6_c74_n34_c)
    );

    fa fa_s6_c75_n35 (
        .a(stage6_col75[0]),
        .b(stage6_col75[1]),
        .c_in(stage6_col75[2]),
        .s(fa_s6_c75_n35_s),
        .c_out(fa_s6_c75_n35_c)
    );

    fa fa_s6_c76_n36 (
        .a(stage6_col76[0]),
        .b(stage6_col76[1]),
        .c_in(stage6_col76[2]),
        .s(fa_s6_c76_n36_s),
        .c_out(fa_s6_c76_n36_c)
    );

    fa fa_s6_c77_n37 (
        .a(stage6_col77[0]),
        .b(stage6_col77[1]),
        .c_in(stage6_col77[2]),
        .s(fa_s6_c77_n37_s),
        .c_out(fa_s6_c77_n37_c)
    );

    fa fa_s6_c78_n38 (
        .a(stage6_col78[0]),
        .b(stage6_col78[1]),
        .c_in(stage6_col78[2]),
        .s(fa_s6_c78_n38_s),
        .c_out(fa_s6_c78_n38_c)
    );

    fa fa_s6_c79_n39 (
        .a(stage6_col79[0]),
        .b(stage6_col79[1]),
        .c_in(stage6_col79[2]),
        .s(fa_s6_c79_n39_s),
        .c_out(fa_s6_c79_n39_c)
    );

    fa fa_s6_c80_n40 (
        .a(stage6_col80[0]),
        .b(stage6_col80[1]),
        .c_in(stage6_col80[2]),
        .s(fa_s6_c80_n40_s),
        .c_out(fa_s6_c80_n40_c)
    );

    fa fa_s6_c81_n41 (
        .a(stage6_col81[0]),
        .b(stage6_col81[1]),
        .c_in(stage6_col81[2]),
        .s(fa_s6_c81_n41_s),
        .c_out(fa_s6_c81_n41_c)
    );

    fa fa_s6_c82_n42 (
        .a(stage6_col82[0]),
        .b(stage6_col82[1]),
        .c_in(stage6_col82[2]),
        .s(fa_s6_c82_n42_s),
        .c_out(fa_s6_c82_n42_c)
    );

    fa fa_s6_c83_n43 (
        .a(stage6_col83[0]),
        .b(stage6_col83[1]),
        .c_in(stage6_col83[2]),
        .s(fa_s6_c83_n43_s),
        .c_out(fa_s6_c83_n43_c)
    );

    fa fa_s6_c84_n44 (
        .a(stage6_col84[0]),
        .b(stage6_col84[1]),
        .c_in(stage6_col84[2]),
        .s(fa_s6_c84_n44_s),
        .c_out(fa_s6_c84_n44_c)
    );

    fa fa_s6_c85_n45 (
        .a(stage6_col85[0]),
        .b(stage6_col85[1]),
        .c_in(stage6_col85[2]),
        .s(fa_s6_c85_n45_s),
        .c_out(fa_s6_c85_n45_c)
    );

    fa fa_s6_c86_n46 (
        .a(stage6_col86[0]),
        .b(stage6_col86[1]),
        .c_in(stage6_col86[2]),
        .s(fa_s6_c86_n46_s),
        .c_out(fa_s6_c86_n46_c)
    );

    fa fa_s6_c87_n47 (
        .a(stage6_col87[0]),
        .b(stage6_col87[1]),
        .c_in(stage6_col87[2]),
        .s(fa_s6_c87_n47_s),
        .c_out(fa_s6_c87_n47_c)
    );

    fa fa_s6_c88_n48 (
        .a(stage6_col88[0]),
        .b(stage6_col88[1]),
        .c_in(stage6_col88[2]),
        .s(fa_s6_c88_n48_s),
        .c_out(fa_s6_c88_n48_c)
    );

    fa fa_s6_c89_n49 (
        .a(stage6_col89[0]),
        .b(stage6_col89[1]),
        .c_in(stage6_col89[2]),
        .s(fa_s6_c89_n49_s),
        .c_out(fa_s6_c89_n49_c)
    );

    fa fa_s6_c90_n50 (
        .a(stage6_col90[0]),
        .b(stage6_col90[1]),
        .c_in(stage6_col90[2]),
        .s(fa_s6_c90_n50_s),
        .c_out(fa_s6_c90_n50_c)
    );

    fa fa_s6_c91_n51 (
        .a(stage6_col91[0]),
        .b(stage6_col91[1]),
        .c_in(stage6_col91[2]),
        .s(fa_s6_c91_n51_s),
        .c_out(fa_s6_c91_n51_c)
    );

    fa fa_s6_c92_n52 (
        .a(stage6_col92[0]),
        .b(stage6_col92[1]),
        .c_in(stage6_col92[2]),
        .s(fa_s6_c92_n52_s),
        .c_out(fa_s6_c92_n52_c)
    );

    fa fa_s6_c93_n53 (
        .a(stage6_col93[0]),
        .b(stage6_col93[1]),
        .c_in(stage6_col93[2]),
        .s(fa_s6_c93_n53_s),
        .c_out(fa_s6_c93_n53_c)
    );

    fa fa_s6_c94_n54 (
        .a(stage6_col94[0]),
        .b(stage6_col94[1]),
        .c_in(stage6_col94[2]),
        .s(fa_s6_c94_n54_s),
        .c_out(fa_s6_c94_n54_c)
    );

    fa fa_s6_c95_n55 (
        .a(stage6_col95[0]),
        .b(stage6_col95[1]),
        .c_in(stage6_col95[2]),
        .s(fa_s6_c95_n55_s),
        .c_out(fa_s6_c95_n55_c)
    );

    fa fa_s6_c96_n56 (
        .a(stage6_col96[0]),
        .b(stage6_col96[1]),
        .c_in(stage6_col96[2]),
        .s(fa_s6_c96_n56_s),
        .c_out(fa_s6_c96_n56_c)
    );

    fa fa_s6_c97_n57 (
        .a(stage6_col97[0]),
        .b(stage6_col97[1]),
        .c_in(stage6_col97[2]),
        .s(fa_s6_c97_n57_s),
        .c_out(fa_s6_c97_n57_c)
    );

    fa fa_s6_c98_n58 (
        .a(stage6_col98[0]),
        .b(stage6_col98[1]),
        .c_in(stage6_col98[2]),
        .s(fa_s6_c98_n58_s),
        .c_out(fa_s6_c98_n58_c)
    );

    fa fa_s6_c99_n59 (
        .a(stage6_col99[0]),
        .b(stage6_col99[1]),
        .c_in(stage6_col99[2]),
        .s(fa_s6_c99_n59_s),
        .c_out(fa_s6_c99_n59_c)
    );

    fa fa_s6_c100_n60 (
        .a(stage6_col100[0]),
        .b(stage6_col100[1]),
        .c_in(stage6_col100[2]),
        .s(fa_s6_c100_n60_s),
        .c_out(fa_s6_c100_n60_c)
    );

    fa fa_s6_c101_n61 (
        .a(stage6_col101[0]),
        .b(stage6_col101[1]),
        .c_in(stage6_col101[2]),
        .s(fa_s6_c101_n61_s),
        .c_out(fa_s6_c101_n61_c)
    );

    fa fa_s6_c102_n62 (
        .a(stage6_col102[0]),
        .b(stage6_col102[1]),
        .c_in(stage6_col102[2]),
        .s(fa_s6_c102_n62_s),
        .c_out(fa_s6_c102_n62_c)
    );

    fa fa_s6_c103_n63 (
        .a(stage6_col103[0]),
        .b(stage6_col103[1]),
        .c_in(stage6_col103[2]),
        .s(fa_s6_c103_n63_s),
        .c_out(fa_s6_c103_n63_c)
    );

    fa fa_s6_c104_n64 (
        .a(stage6_col104[0]),
        .b(stage6_col104[1]),
        .c_in(stage6_col104[2]),
        .s(fa_s6_c104_n64_s),
        .c_out(fa_s6_c104_n64_c)
    );

    fa fa_s6_c105_n65 (
        .a(stage6_col105[0]),
        .b(stage6_col105[1]),
        .c_in(stage6_col105[2]),
        .s(fa_s6_c105_n65_s),
        .c_out(fa_s6_c105_n65_c)
    );

    fa fa_s6_c106_n66 (
        .a(stage6_col106[0]),
        .b(stage6_col106[1]),
        .c_in(stage6_col106[2]),
        .s(fa_s6_c106_n66_s),
        .c_out(fa_s6_c106_n66_c)
    );

    fa fa_s6_c107_n67 (
        .a(stage6_col107[0]),
        .b(stage6_col107[1]),
        .c_in(stage6_col107[2]),
        .s(fa_s6_c107_n67_s),
        .c_out(fa_s6_c107_n67_c)
    );

    fa fa_s6_c108_n68 (
        .a(stage6_col108[0]),
        .b(stage6_col108[1]),
        .c_in(stage6_col108[2]),
        .s(fa_s6_c108_n68_s),
        .c_out(fa_s6_c108_n68_c)
    );

    fa fa_s6_c109_n69 (
        .a(stage6_col109[0]),
        .b(stage6_col109[1]),
        .c_in(stage6_col109[2]),
        .s(fa_s6_c109_n69_s),
        .c_out(fa_s6_c109_n69_c)
    );

    fa fa_s6_c110_n70 (
        .a(stage6_col110[0]),
        .b(stage6_col110[1]),
        .c_in(stage6_col110[2]),
        .s(fa_s6_c110_n70_s),
        .c_out(fa_s6_c110_n70_c)
    );

    fa fa_s6_c111_n71 (
        .a(stage6_col111[0]),
        .b(stage6_col111[1]),
        .c_in(stage6_col111[2]),
        .s(fa_s6_c111_n71_s),
        .c_out(fa_s6_c111_n71_c)
    );

    fa fa_s6_c112_n72 (
        .a(stage6_col112[0]),
        .b(stage6_col112[1]),
        .c_in(stage6_col112[2]),
        .s(fa_s6_c112_n72_s),
        .c_out(fa_s6_c112_n72_c)
    );

    fa fa_s6_c113_n73 (
        .a(stage6_col113[0]),
        .b(stage6_col113[1]),
        .c_in(stage6_col113[2]),
        .s(fa_s6_c113_n73_s),
        .c_out(fa_s6_c113_n73_c)
    );

    fa fa_s6_c114_n74 (
        .a(stage6_col114[0]),
        .b(stage6_col114[1]),
        .c_in(stage6_col114[2]),
        .s(fa_s6_c114_n74_s),
        .c_out(fa_s6_c114_n74_c)
    );

    fa fa_s6_c115_n75 (
        .a(stage6_col115[0]),
        .b(stage6_col115[1]),
        .c_in(stage6_col115[2]),
        .s(fa_s6_c115_n75_s),
        .c_out(fa_s6_c115_n75_c)
    );

    fa fa_s6_c116_n76 (
        .a(stage6_col116[0]),
        .b(stage6_col116[1]),
        .c_in(stage6_col116[2]),
        .s(fa_s6_c116_n76_s),
        .c_out(fa_s6_c116_n76_c)
    );

    fa fa_s6_c117_n77 (
        .a(stage6_col117[0]),
        .b(stage6_col117[1]),
        .c_in(stage6_col117[2]),
        .s(fa_s6_c117_n77_s),
        .c_out(fa_s6_c117_n77_c)
    );

    fa fa_s6_c118_n78 (
        .a(stage6_col118[0]),
        .b(stage6_col118[1]),
        .c_in(stage6_col118[2]),
        .s(fa_s6_c118_n78_s),
        .c_out(fa_s6_c118_n78_c)
    );

    fa fa_s6_c119_n79 (
        .a(stage6_col119[0]),
        .b(stage6_col119[1]),
        .c_in(stage6_col119[2]),
        .s(fa_s6_c119_n79_s),
        .c_out(fa_s6_c119_n79_c)
    );

    fa fa_s6_c120_n80 (
        .a(stage6_col120[0]),
        .b(stage6_col120[1]),
        .c_in(stage6_col120[2]),
        .s(fa_s6_c120_n80_s),
        .c_out(fa_s6_c120_n80_c)
    );

    fa fa_s6_c121_n81 (
        .a(stage6_col121[0]),
        .b(stage6_col121[1]),
        .c_in(stage6_col121[2]),
        .s(fa_s6_c121_n81_s),
        .c_out(fa_s6_c121_n81_c)
    );

    fa fa_s6_c122_n82 (
        .a(stage6_col122[0]),
        .b(stage6_col122[1]),
        .c_in(stage6_col122[2]),
        .s(fa_s6_c122_n82_s),
        .c_out(fa_s6_c122_n82_c)
    );

    fa fa_s6_c123_n83 (
        .a(stage6_col123[0]),
        .b(stage6_col123[1]),
        .c_in(stage6_col123[2]),
        .s(fa_s6_c123_n83_s),
        .c_out(fa_s6_c123_n83_c)
    );

    fa fa_s6_c124_n84 (
        .a(stage6_col124[0]),
        .b(stage6_col124[1]),
        .c_in(stage6_col124[2]),
        .s(fa_s6_c124_n84_s),
        .c_out(fa_s6_c124_n84_c)
    );

    fa fa_s6_c125_n85 (
        .a(stage6_col125[0]),
        .b(stage6_col125[1]),
        .c_in(stage6_col125[2]),
        .s(fa_s6_c125_n85_s),
        .c_out(fa_s6_c125_n85_c)
    );

    fa fa_s6_c126_n86 (
        .a(stage6_col126[0]),
        .b(stage6_col126[1]),
        .c_in(stage6_col126[2]),
        .s(fa_s6_c126_n86_s),
        .c_out(fa_s6_c126_n86_c)
    );

    ha ha_s6_c6_n0 (
        .a(stage6_col6[0]),
        .b(stage6_col6[1]),
        .s(ha_s6_c6_n0_s),
        .c_out(ha_s6_c6_n0_c)
    );

    // Map to Stage 7 columns
    generate
        if (PIPE) begin : gen_stage7_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage7_col0[0] <= 1'b0;
                    stage7_col1[0] <= 1'b0;
                    stage7_col2[0] <= 1'b0;
                    stage7_col3[0] <= 1'b0;
                    stage7_col4[0] <= 1'b0;
                    stage7_col5[0] <= 1'b0;
                    stage7_col6[0] <= 1'b0;
                    stage7_col7[0] <= 1'b0;
                    stage7_col7[1] <= 1'b0;
                    stage7_col8[0] <= 1'b0;
                    stage7_col9[0] <= 1'b0;
                    stage7_col9[1] <= 1'b0;
                    stage7_col9[2] <= 1'b0;
                    stage7_col10[0] <= 1'b0;
                    stage7_col10[1] <= 1'b0;
                    stage7_col11[0] <= 1'b0;
                    stage7_col11[1] <= 1'b0;
                    stage7_col12[0] <= 1'b0;
                    stage7_col12[1] <= 1'b0;
                    stage7_col13[0] <= 1'b0;
                    stage7_col13[1] <= 1'b0;
                    stage7_col14[0] <= 1'b0;
                    stage7_col14[1] <= 1'b0;
                    stage7_col15[0] <= 1'b0;
                    stage7_col15[1] <= 1'b0;
                    stage7_col16[0] <= 1'b0;
                    stage7_col16[1] <= 1'b0;
                    stage7_col17[0] <= 1'b0;
                    stage7_col17[1] <= 1'b0;
                    stage7_col18[0] <= 1'b0;
                    stage7_col18[1] <= 1'b0;
                    stage7_col19[0] <= 1'b0;
                    stage7_col19[1] <= 1'b0;
                    stage7_col20[0] <= 1'b0;
                    stage7_col20[1] <= 1'b0;
                    stage7_col21[0] <= 1'b0;
                    stage7_col21[1] <= 1'b0;
                    stage7_col22[0] <= 1'b0;
                    stage7_col22[1] <= 1'b0;
                    stage7_col23[0] <= 1'b0;
                    stage7_col23[1] <= 1'b0;
                    stage7_col24[0] <= 1'b0;
                    stage7_col24[1] <= 1'b0;
                    stage7_col25[0] <= 1'b0;
                    stage7_col25[1] <= 1'b0;
                    stage7_col26[0] <= 1'b0;
                    stage7_col26[1] <= 1'b0;
                    stage7_col27[0] <= 1'b0;
                    stage7_col27[1] <= 1'b0;
                    stage7_col28[0] <= 1'b0;
                    stage7_col28[1] <= 1'b0;
                    stage7_col29[0] <= 1'b0;
                    stage7_col29[1] <= 1'b0;
                    stage7_col30[0] <= 1'b0;
                    stage7_col30[1] <= 1'b0;
                    stage7_col31[0] <= 1'b0;
                    stage7_col31[1] <= 1'b0;
                    stage7_col32[0] <= 1'b0;
                    stage7_col32[1] <= 1'b0;
                    stage7_col33[0] <= 1'b0;
                    stage7_col33[1] <= 1'b0;
                    stage7_col34[0] <= 1'b0;
                    stage7_col34[1] <= 1'b0;
                    stage7_col35[0] <= 1'b0;
                    stage7_col35[1] <= 1'b0;
                    stage7_col36[0] <= 1'b0;
                    stage7_col36[1] <= 1'b0;
                    stage7_col37[0] <= 1'b0;
                    stage7_col37[1] <= 1'b0;
                    stage7_col38[0] <= 1'b0;
                    stage7_col38[1] <= 1'b0;
                    stage7_col39[0] <= 1'b0;
                    stage7_col39[1] <= 1'b0;
                    stage7_col40[0] <= 1'b0;
                    stage7_col40[1] <= 1'b0;
                    stage7_col41[0] <= 1'b0;
                    stage7_col41[1] <= 1'b0;
                    stage7_col42[0] <= 1'b0;
                    stage7_col42[1] <= 1'b0;
                    stage7_col43[0] <= 1'b0;
                    stage7_col43[1] <= 1'b0;
                    stage7_col44[0] <= 1'b0;
                    stage7_col44[1] <= 1'b0;
                    stage7_col45[0] <= 1'b0;
                    stage7_col45[1] <= 1'b0;
                    stage7_col46[0] <= 1'b0;
                    stage7_col46[1] <= 1'b0;
                    stage7_col47[0] <= 1'b0;
                    stage7_col47[1] <= 1'b0;
                    stage7_col48[0] <= 1'b0;
                    stage7_col48[1] <= 1'b0;
                    stage7_col49[0] <= 1'b0;
                    stage7_col49[1] <= 1'b0;
                    stage7_col50[0] <= 1'b0;
                    stage7_col50[1] <= 1'b0;
                    stage7_col51[0] <= 1'b0;
                    stage7_col51[1] <= 1'b0;
                    stage7_col52[0] <= 1'b0;
                    stage7_col52[1] <= 1'b0;
                    stage7_col53[0] <= 1'b0;
                    stage7_col53[1] <= 1'b0;
                    stage7_col54[0] <= 1'b0;
                    stage7_col54[1] <= 1'b0;
                    stage7_col55[0] <= 1'b0;
                    stage7_col55[1] <= 1'b0;
                    stage7_col56[0] <= 1'b0;
                    stage7_col56[1] <= 1'b0;
                    stage7_col57[0] <= 1'b0;
                    stage7_col57[1] <= 1'b0;
                    stage7_col58[0] <= 1'b0;
                    stage7_col58[1] <= 1'b0;
                    stage7_col59[0] <= 1'b0;
                    stage7_col59[1] <= 1'b0;
                    stage7_col60[0] <= 1'b0;
                    stage7_col60[1] <= 1'b0;
                    stage7_col60[2] <= 1'b0;
                    stage7_col61[0] <= 1'b0;
                    stage7_col61[1] <= 1'b0;
                    stage7_col61[2] <= 1'b0;
                    stage7_col62[0] <= 1'b0;
                    stage7_col62[1] <= 1'b0;
                    stage7_col62[2] <= 1'b0;
                    stage7_col63[0] <= 1'b0;
                    stage7_col63[1] <= 1'b0;
                    stage7_col63[2] <= 1'b0;
                    stage7_col64[0] <= 1'b0;
                    stage7_col64[1] <= 1'b0;
                    stage7_col64[2] <= 1'b0;
                    stage7_col65[0] <= 1'b0;
                    stage7_col65[1] <= 1'b0;
                    stage7_col65[2] <= 1'b0;
                    stage7_col66[0] <= 1'b0;
                    stage7_col66[1] <= 1'b0;
                    stage7_col66[2] <= 1'b0;
                    stage7_col67[0] <= 1'b0;
                    stage7_col67[1] <= 1'b0;
                    stage7_col67[2] <= 1'b0;
                    stage7_col68[0] <= 1'b0;
                    stage7_col68[1] <= 1'b0;
                    stage7_col68[2] <= 1'b0;
                    stage7_col69[0] <= 1'b0;
                    stage7_col69[1] <= 1'b0;
                    stage7_col69[2] <= 1'b0;
                    stage7_col70[0] <= 1'b0;
                    stage7_col70[1] <= 1'b0;
                    stage7_col70[2] <= 1'b0;
                    stage7_col71[0] <= 1'b0;
                    stage7_col71[1] <= 1'b0;
                    stage7_col71[2] <= 1'b0;
                    stage7_col72[0] <= 1'b0;
                    stage7_col72[1] <= 1'b0;
                    stage7_col72[2] <= 1'b0;
                    stage7_col73[0] <= 1'b0;
                    stage7_col73[1] <= 1'b0;
                    stage7_col73[2] <= 1'b0;
                    stage7_col74[0] <= 1'b0;
                    stage7_col74[1] <= 1'b0;
                    stage7_col74[2] <= 1'b0;
                    stage7_col75[0] <= 1'b0;
                    stage7_col75[1] <= 1'b0;
                    stage7_col75[2] <= 1'b0;
                    stage7_col76[0] <= 1'b0;
                    stage7_col76[1] <= 1'b0;
                    stage7_col76[2] <= 1'b0;
                    stage7_col77[0] <= 1'b0;
                    stage7_col77[1] <= 1'b0;
                    stage7_col77[2] <= 1'b0;
                    stage7_col78[0] <= 1'b0;
                    stage7_col78[1] <= 1'b0;
                    stage7_col78[2] <= 1'b0;
                    stage7_col79[0] <= 1'b0;
                    stage7_col79[1] <= 1'b0;
                    stage7_col79[2] <= 1'b0;
                    stage7_col80[0] <= 1'b0;
                    stage7_col80[1] <= 1'b0;
                    stage7_col80[2] <= 1'b0;
                    stage7_col81[0] <= 1'b0;
                    stage7_col81[1] <= 1'b0;
                    stage7_col81[2] <= 1'b0;
                    stage7_col82[0] <= 1'b0;
                    stage7_col82[1] <= 1'b0;
                    stage7_col82[2] <= 1'b0;
                    stage7_col83[0] <= 1'b0;
                    stage7_col83[1] <= 1'b0;
                    stage7_col83[2] <= 1'b0;
                    stage7_col84[0] <= 1'b0;
                    stage7_col84[1] <= 1'b0;
                    stage7_col84[2] <= 1'b0;
                    stage7_col85[0] <= 1'b0;
                    stage7_col85[1] <= 1'b0;
                    stage7_col85[2] <= 1'b0;
                    stage7_col86[0] <= 1'b0;
                    stage7_col86[1] <= 1'b0;
                    stage7_col86[2] <= 1'b0;
                    stage7_col87[0] <= 1'b0;
                    stage7_col87[1] <= 1'b0;
                    stage7_col87[2] <= 1'b0;
                    stage7_col88[0] <= 1'b0;
                    stage7_col88[1] <= 1'b0;
                    stage7_col88[2] <= 1'b0;
                    stage7_col89[0] <= 1'b0;
                    stage7_col89[1] <= 1'b0;
                    stage7_col89[2] <= 1'b0;
                    stage7_col90[0] <= 1'b0;
                    stage7_col90[1] <= 1'b0;
                    stage7_col90[2] <= 1'b0;
                    stage7_col91[0] <= 1'b0;
                    stage7_col91[1] <= 1'b0;
                    stage7_col91[2] <= 1'b0;
                    stage7_col92[0] <= 1'b0;
                    stage7_col92[1] <= 1'b0;
                    stage7_col92[2] <= 1'b0;
                    stage7_col93[0] <= 1'b0;
                    stage7_col93[1] <= 1'b0;
                    stage7_col93[2] <= 1'b0;
                    stage7_col94[0] <= 1'b0;
                    stage7_col94[1] <= 1'b0;
                    stage7_col94[2] <= 1'b0;
                    stage7_col95[0] <= 1'b0;
                    stage7_col95[1] <= 1'b0;
                    stage7_col95[2] <= 1'b0;
                    stage7_col96[0] <= 1'b0;
                    stage7_col96[1] <= 1'b0;
                    stage7_col96[2] <= 1'b0;
                    stage7_col97[0] <= 1'b0;
                    stage7_col97[1] <= 1'b0;
                    stage7_col97[2] <= 1'b0;
                    stage7_col98[0] <= 1'b0;
                    stage7_col98[1] <= 1'b0;
                    stage7_col98[2] <= 1'b0;
                    stage7_col99[0] <= 1'b0;
                    stage7_col99[1] <= 1'b0;
                    stage7_col99[2] <= 1'b0;
                    stage7_col100[0] <= 1'b0;
                    stage7_col100[1] <= 1'b0;
                    stage7_col100[2] <= 1'b0;
                    stage7_col101[0] <= 1'b0;
                    stage7_col101[1] <= 1'b0;
                    stage7_col101[2] <= 1'b0;
                    stage7_col102[0] <= 1'b0;
                    stage7_col102[1] <= 1'b0;
                    stage7_col102[2] <= 1'b0;
                    stage7_col103[0] <= 1'b0;
                    stage7_col103[1] <= 1'b0;
                    stage7_col103[2] <= 1'b0;
                    stage7_col104[0] <= 1'b0;
                    stage7_col104[1] <= 1'b0;
                    stage7_col104[2] <= 1'b0;
                    stage7_col105[0] <= 1'b0;
                    stage7_col105[1] <= 1'b0;
                    stage7_col105[2] <= 1'b0;
                    stage7_col106[0] <= 1'b0;
                    stage7_col106[1] <= 1'b0;
                    stage7_col106[2] <= 1'b0;
                    stage7_col107[0] <= 1'b0;
                    stage7_col107[1] <= 1'b0;
                    stage7_col107[2] <= 1'b0;
                    stage7_col108[0] <= 1'b0;
                    stage7_col108[1] <= 1'b0;
                    stage7_col108[2] <= 1'b0;
                    stage7_col109[0] <= 1'b0;
                    stage7_col109[1] <= 1'b0;
                    stage7_col109[2] <= 1'b0;
                    stage7_col110[0] <= 1'b0;
                    stage7_col110[1] <= 1'b0;
                    stage7_col110[2] <= 1'b0;
                    stage7_col111[0] <= 1'b0;
                    stage7_col111[1] <= 1'b0;
                    stage7_col111[2] <= 1'b0;
                    stage7_col112[0] <= 1'b0;
                    stage7_col112[1] <= 1'b0;
                    stage7_col112[2] <= 1'b0;
                    stage7_col113[0] <= 1'b0;
                    stage7_col113[1] <= 1'b0;
                    stage7_col113[2] <= 1'b0;
                    stage7_col114[0] <= 1'b0;
                    stage7_col114[1] <= 1'b0;
                    stage7_col114[2] <= 1'b0;
                    stage7_col115[0] <= 1'b0;
                    stage7_col115[1] <= 1'b0;
                    stage7_col115[2] <= 1'b0;
                    stage7_col116[0] <= 1'b0;
                    stage7_col116[1] <= 1'b0;
                    stage7_col116[2] <= 1'b0;
                    stage7_col117[0] <= 1'b0;
                    stage7_col117[1] <= 1'b0;
                    stage7_col117[2] <= 1'b0;
                    stage7_col118[0] <= 1'b0;
                    stage7_col118[1] <= 1'b0;
                    stage7_col118[2] <= 1'b0;
                    stage7_col119[0] <= 1'b0;
                    stage7_col119[1] <= 1'b0;
                    stage7_col119[2] <= 1'b0;
                    stage7_col120[0] <= 1'b0;
                    stage7_col120[1] <= 1'b0;
                    stage7_col120[2] <= 1'b0;
                    stage7_col121[0] <= 1'b0;
                    stage7_col121[1] <= 1'b0;
                    stage7_col121[2] <= 1'b0;
                    stage7_col122[0] <= 1'b0;
                    stage7_col122[1] <= 1'b0;
                    stage7_col122[2] <= 1'b0;
                    stage7_col123[0] <= 1'b0;
                    stage7_col123[1] <= 1'b0;
                    stage7_col123[2] <= 1'b0;
                    stage7_col124[0] <= 1'b0;
                    stage7_col124[1] <= 1'b0;
                    stage7_col124[2] <= 1'b0;
                    stage7_col125[0] <= 1'b0;
                    stage7_col125[1] <= 1'b0;
                    stage7_col125[2] <= 1'b0;
                    stage7_col126[0] <= 1'b0;
                    stage7_col126[1] <= 1'b0;
                    stage7_col126[2] <= 1'b0;
                    stage7_col127[0] <= 1'b0;
                    stage7_col127[1] <= 1'b0;
                    stage7_col127[2] <= 1'b0;
                    stage7_col127[3] <= 1'b0;
                    stage7_col127[4] <= 1'b0;
                    stage7_col127[5] <= 1'b0;
                    stage7_col127[6] <= 1'b0;
                    stage7_col127[7] <= 1'b0;
                    stage7_col127[8] <= 1'b0;
                    stage7_col127[9] <= 1'b0;
                    stage7_col127[10] <= 1'b0;
                    stage7_col127[11] <= 1'b0;
                    stage7_col127[12] <= 1'b0;
                    stage7_col127[13] <= 1'b0;
                    stage7_col127[14] <= 1'b0;
                    stage7_col127[15] <= 1'b0;
                    stage7_col127[16] <= 1'b0;
                    stage7_col127[17] <= 1'b0;
                    stage7_col127[18] <= 1'b0;
                    stage7_col127[19] <= 1'b0;
                    stage7_col127[20] <= 1'b0;
                    stage7_col127[21] <= 1'b0;
                    stage7_col127[22] <= 1'b0;
                    stage7_col127[23] <= 1'b0;
                    stage7_col127[24] <= 1'b0;
                    stage7_col127[25] <= 1'b0;
                    stage7_col127[26] <= 1'b0;
                    stage7_col127[27] <= 1'b0;
                    stage7_col127[28] <= 1'b0;
                    stage7_col127[29] <= 1'b0;
                    stage7_col127[30] <= 1'b0;
                    stage7_col127[31] <= 1'b0;
                    stage7_col127[32] <= 1'b0;
                    stage7_col127[33] <= 1'b0;
                    stage7_col127[34] <= 1'b0;
                    stage7_col127[35] <= 1'b0;
                    stage7_col127[36] <= 1'b0;
                    stage7_col127[37] <= 1'b0;
                    stage7_col127[38] <= 1'b0;
                    stage7_col127[39] <= 1'b0;
                    stage7_col127[40] <= 1'b0;
                    stage7_col127[41] <= 1'b0;
                    stage7_col127[42] <= 1'b0;
                    stage7_col127[43] <= 1'b0;
                    stage7_col127[44] <= 1'b0;
                    stage7_col127[45] <= 1'b0;
                    stage7_col127[46] <= 1'b0;
                    stage7_col127[47] <= 1'b0;
                    stage7_col127[48] <= 1'b0;
                    stage7_col127[49] <= 1'b0;
                    stage7_col127[50] <= 1'b0;
                    stage7_col127[51] <= 1'b0;
                    stage7_col127[52] <= 1'b0;
                    stage7_col127[53] <= 1'b0;
                    stage7_col127[54] <= 1'b0;
                    stage7_col127[55] <= 1'b0;
                    stage7_col127[56] <= 1'b0;
                    stage7_col127[57] <= 1'b0;
                    stage7_col127[58] <= 1'b0;
                    stage7_col127[59] <= 1'b0;
                    stage7_col127[60] <= 1'b0;
                    stage7_col127[61] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage7_col0[0] <= stage6_col0[0];
                    stage7_col1[0] <= stage6_col1[0];
                    stage7_col2[0] <= stage6_col2[0];
                    stage7_col3[0] <= stage6_col3[0];
                    stage7_col4[0] <= stage6_col4[0];
                    stage7_col5[0] <= stage6_col5[0];
                    stage7_col6[0] <= ha_s6_c6_n0_s;
                    stage7_col7[0] <= ha_s6_c6_n0_c;
                    stage7_col7[1] <= stage6_col7[0];
                    stage7_col8[0] <= fa_s6_c8_n0_s;
                    stage7_col9[0] <= fa_s6_c8_n0_c;
                    stage7_col9[1] <= stage6_col9[0];
                    stage7_col9[2] <= stage6_col9[1];
                    stage7_col10[0] <= stage6_col10[0];
                    stage7_col10[1] <= stage6_col10[1];
                    stage7_col11[0] <= stage6_col11[0];
                    stage7_col11[1] <= stage6_col11[1];
                    stage7_col12[0] <= stage6_col12[0];
                    stage7_col12[1] <= stage6_col12[1];
                    stage7_col13[0] <= stage6_col13[0];
                    stage7_col13[1] <= stage6_col13[1];
                    stage7_col14[0] <= stage6_col14[0];
                    stage7_col14[1] <= stage6_col14[1];
                    stage7_col15[0] <= stage6_col15[0];
                    stage7_col15[1] <= stage6_col15[1];
                    stage7_col16[0] <= stage6_col16[0];
                    stage7_col16[1] <= stage6_col16[1];
                    stage7_col17[0] <= stage6_col17[0];
                    stage7_col17[1] <= stage6_col17[1];
                    stage7_col18[0] <= stage6_col18[0];
                    stage7_col18[1] <= stage6_col18[1];
                    stage7_col19[0] <= stage6_col19[0];
                    stage7_col19[1] <= stage6_col19[1];
                    stage7_col20[0] <= stage6_col20[0];
                    stage7_col20[1] <= stage6_col20[1];
                    stage7_col21[0] <= stage6_col21[0];
                    stage7_col21[1] <= stage6_col21[1];
                    stage7_col22[0] <= stage6_col22[0];
                    stage7_col22[1] <= stage6_col22[1];
                    stage7_col23[0] <= stage6_col23[0];
                    stage7_col23[1] <= stage6_col23[1];
                    stage7_col24[0] <= stage6_col24[0];
                    stage7_col24[1] <= stage6_col24[1];
                    stage7_col25[0] <= stage6_col25[0];
                    stage7_col25[1] <= stage6_col25[1];
                    stage7_col26[0] <= stage6_col26[0];
                    stage7_col26[1] <= stage6_col26[1];
                    stage7_col27[0] <= stage6_col27[0];
                    stage7_col27[1] <= stage6_col27[1];
                    stage7_col28[0] <= stage6_col28[0];
                    stage7_col28[1] <= stage6_col28[1];
                    stage7_col29[0] <= stage6_col29[0];
                    stage7_col29[1] <= stage6_col29[1];
                    stage7_col30[0] <= stage6_col30[0];
                    stage7_col30[1] <= stage6_col30[1];
                    stage7_col31[0] <= stage6_col31[0];
                    stage7_col31[1] <= stage6_col31[1];
                    stage7_col32[0] <= stage6_col32[0];
                    stage7_col32[1] <= stage6_col32[1];
                    stage7_col33[0] <= stage6_col33[0];
                    stage7_col33[1] <= stage6_col33[1];
                    stage7_col34[0] <= stage6_col34[0];
                    stage7_col34[1] <= stage6_col34[1];
                    stage7_col35[0] <= stage6_col35[0];
                    stage7_col35[1] <= stage6_col35[1];
                    stage7_col36[0] <= stage6_col36[0];
                    stage7_col36[1] <= stage6_col36[1];
                    stage7_col37[0] <= stage6_col37[0];
                    stage7_col37[1] <= stage6_col37[1];
                    stage7_col38[0] <= stage6_col38[0];
                    stage7_col38[1] <= stage6_col38[1];
                    stage7_col39[0] <= stage6_col39[0];
                    stage7_col39[1] <= stage6_col39[1];
                    stage7_col40[0] <= stage6_col40[0];
                    stage7_col40[1] <= stage6_col40[1];
                    stage7_col41[0] <= fa_s6_c41_n1_s;
                    stage7_col41[1] <= stage6_col41[3];
                    stage7_col42[0] <= fa_s6_c41_n1_c;
                    stage7_col42[1] <= fa_s6_c42_n2_s;
                    stage7_col43[0] <= fa_s6_c42_n2_c;
                    stage7_col43[1] <= fa_s6_c43_n3_s;
                    stage7_col44[0] <= fa_s6_c43_n3_c;
                    stage7_col44[1] <= fa_s6_c44_n4_s;
                    stage7_col45[0] <= fa_s6_c44_n4_c;
                    stage7_col45[1] <= fa_s6_c45_n5_s;
                    stage7_col46[0] <= fa_s6_c45_n5_c;
                    stage7_col46[1] <= fa_s6_c46_n6_s;
                    stage7_col47[0] <= fa_s6_c46_n6_c;
                    stage7_col47[1] <= fa_s6_c47_n7_s;
                    stage7_col48[0] <= fa_s6_c47_n7_c;
                    stage7_col48[1] <= fa_s6_c48_n8_s;
                    stage7_col49[0] <= fa_s6_c48_n8_c;
                    stage7_col49[1] <= fa_s6_c49_n9_s;
                    stage7_col50[0] <= fa_s6_c49_n9_c;
                    stage7_col50[1] <= fa_s6_c50_n10_s;
                    stage7_col51[0] <= fa_s6_c50_n10_c;
                    stage7_col51[1] <= fa_s6_c51_n11_s;
                    stage7_col52[0] <= fa_s6_c51_n11_c;
                    stage7_col52[1] <= fa_s6_c52_n12_s;
                    stage7_col53[0] <= fa_s6_c52_n12_c;
                    stage7_col53[1] <= fa_s6_c53_n13_s;
                    stage7_col54[0] <= fa_s6_c53_n13_c;
                    stage7_col54[1] <= fa_s6_c54_n14_s;
                    stage7_col55[0] <= fa_s6_c54_n14_c;
                    stage7_col55[1] <= fa_s6_c55_n15_s;
                    stage7_col56[0] <= fa_s6_c55_n15_c;
                    stage7_col56[1] <= fa_s6_c56_n16_s;
                    stage7_col57[0] <= fa_s6_c56_n16_c;
                    stage7_col57[1] <= fa_s6_c57_n17_s;
                    stage7_col58[0] <= fa_s6_c57_n17_c;
                    stage7_col58[1] <= fa_s6_c58_n18_s;
                    stage7_col59[0] <= fa_s6_c58_n18_c;
                    stage7_col59[1] <= fa_s6_c59_n19_s;
                    stage7_col60[0] <= fa_s6_c59_n19_c;
                    stage7_col60[1] <= fa_s6_c60_n20_s;
                    stage7_col60[2] <= stage6_col60[3];
                    stage7_col61[0] <= fa_s6_c60_n20_c;
                    stage7_col61[1] <= fa_s6_c61_n21_s;
                    stage7_col61[2] <= stage6_col61[3];
                    stage7_col62[0] <= fa_s6_c61_n21_c;
                    stage7_col62[1] <= fa_s6_c62_n22_s;
                    stage7_col62[2] <= stage6_col62[3];
                    stage7_col63[0] <= fa_s6_c62_n22_c;
                    stage7_col63[1] <= fa_s6_c63_n23_s;
                    stage7_col63[2] <= stage6_col63[3];
                    stage7_col64[0] <= fa_s6_c63_n23_c;
                    stage7_col64[1] <= fa_s6_c64_n24_s;
                    stage7_col64[2] <= stage6_col64[3];
                    stage7_col65[0] <= fa_s6_c64_n24_c;
                    stage7_col65[1] <= fa_s6_c65_n25_s;
                    stage7_col65[2] <= stage6_col65[3];
                    stage7_col66[0] <= fa_s6_c65_n25_c;
                    stage7_col66[1] <= fa_s6_c66_n26_s;
                    stage7_col66[2] <= stage6_col66[3];
                    stage7_col67[0] <= fa_s6_c66_n26_c;
                    stage7_col67[1] <= fa_s6_c67_n27_s;
                    stage7_col67[2] <= stage6_col67[3];
                    stage7_col68[0] <= fa_s6_c67_n27_c;
                    stage7_col68[1] <= fa_s6_c68_n28_s;
                    stage7_col68[2] <= stage6_col68[3];
                    stage7_col69[0] <= fa_s6_c68_n28_c;
                    stage7_col69[1] <= fa_s6_c69_n29_s;
                    stage7_col69[2] <= stage6_col69[3];
                    stage7_col70[0] <= fa_s6_c69_n29_c;
                    stage7_col70[1] <= fa_s6_c70_n30_s;
                    stage7_col70[2] <= stage6_col70[3];
                    stage7_col71[0] <= fa_s6_c70_n30_c;
                    stage7_col71[1] <= fa_s6_c71_n31_s;
                    stage7_col71[2] <= stage6_col71[3];
                    stage7_col72[0] <= fa_s6_c71_n31_c;
                    stage7_col72[1] <= fa_s6_c72_n32_s;
                    stage7_col72[2] <= stage6_col72[3];
                    stage7_col73[0] <= fa_s6_c72_n32_c;
                    stage7_col73[1] <= fa_s6_c73_n33_s;
                    stage7_col73[2] <= stage6_col73[3];
                    stage7_col74[0] <= fa_s6_c73_n33_c;
                    stage7_col74[1] <= fa_s6_c74_n34_s;
                    stage7_col74[2] <= stage6_col74[3];
                    stage7_col75[0] <= fa_s6_c74_n34_c;
                    stage7_col75[1] <= fa_s6_c75_n35_s;
                    stage7_col75[2] <= stage6_col75[3];
                    stage7_col76[0] <= fa_s6_c75_n35_c;
                    stage7_col76[1] <= fa_s6_c76_n36_s;
                    stage7_col76[2] <= stage6_col76[3];
                    stage7_col77[0] <= fa_s6_c76_n36_c;
                    stage7_col77[1] <= fa_s6_c77_n37_s;
                    stage7_col77[2] <= stage6_col77[3];
                    stage7_col78[0] <= fa_s6_c77_n37_c;
                    stage7_col78[1] <= fa_s6_c78_n38_s;
                    stage7_col78[2] <= stage6_col78[3];
                    stage7_col79[0] <= fa_s6_c78_n38_c;
                    stage7_col79[1] <= fa_s6_c79_n39_s;
                    stage7_col79[2] <= stage6_col79[3];
                    stage7_col80[0] <= fa_s6_c79_n39_c;
                    stage7_col80[1] <= fa_s6_c80_n40_s;
                    stage7_col80[2] <= stage6_col80[3];
                    stage7_col81[0] <= fa_s6_c80_n40_c;
                    stage7_col81[1] <= fa_s6_c81_n41_s;
                    stage7_col81[2] <= stage6_col81[3];
                    stage7_col82[0] <= fa_s6_c81_n41_c;
                    stage7_col82[1] <= fa_s6_c82_n42_s;
                    stage7_col82[2] <= stage6_col82[3];
                    stage7_col83[0] <= fa_s6_c82_n42_c;
                    stage7_col83[1] <= fa_s6_c83_n43_s;
                    stage7_col83[2] <= stage6_col83[3];
                    stage7_col84[0] <= fa_s6_c83_n43_c;
                    stage7_col84[1] <= fa_s6_c84_n44_s;
                    stage7_col84[2] <= stage6_col84[3];
                    stage7_col85[0] <= fa_s6_c84_n44_c;
                    stage7_col85[1] <= fa_s6_c85_n45_s;
                    stage7_col85[2] <= stage6_col85[3];
                    stage7_col86[0] <= fa_s6_c85_n45_c;
                    stage7_col86[1] <= fa_s6_c86_n46_s;
                    stage7_col86[2] <= stage6_col86[3];
                    stage7_col87[0] <= fa_s6_c86_n46_c;
                    stage7_col87[1] <= fa_s6_c87_n47_s;
                    stage7_col87[2] <= stage6_col87[3];
                    stage7_col88[0] <= fa_s6_c87_n47_c;
                    stage7_col88[1] <= fa_s6_c88_n48_s;
                    stage7_col88[2] <= stage6_col88[3];
                    stage7_col89[0] <= fa_s6_c88_n48_c;
                    stage7_col89[1] <= fa_s6_c89_n49_s;
                    stage7_col89[2] <= stage6_col89[3];
                    stage7_col90[0] <= fa_s6_c89_n49_c;
                    stage7_col90[1] <= fa_s6_c90_n50_s;
                    stage7_col90[2] <= stage6_col90[3];
                    stage7_col91[0] <= fa_s6_c90_n50_c;
                    stage7_col91[1] <= fa_s6_c91_n51_s;
                    stage7_col91[2] <= stage6_col91[3];
                    stage7_col92[0] <= fa_s6_c91_n51_c;
                    stage7_col92[1] <= fa_s6_c92_n52_s;
                    stage7_col92[2] <= stage6_col92[3];
                    stage7_col93[0] <= fa_s6_c92_n52_c;
                    stage7_col93[1] <= fa_s6_c93_n53_s;
                    stage7_col93[2] <= stage6_col93[3];
                    stage7_col94[0] <= fa_s6_c93_n53_c;
                    stage7_col94[1] <= fa_s6_c94_n54_s;
                    stage7_col94[2] <= stage6_col94[3];
                    stage7_col95[0] <= fa_s6_c94_n54_c;
                    stage7_col95[1] <= fa_s6_c95_n55_s;
                    stage7_col95[2] <= stage6_col95[3];
                    stage7_col96[0] <= fa_s6_c95_n55_c;
                    stage7_col96[1] <= fa_s6_c96_n56_s;
                    stage7_col96[2] <= stage6_col96[3];
                    stage7_col97[0] <= fa_s6_c96_n56_c;
                    stage7_col97[1] <= fa_s6_c97_n57_s;
                    stage7_col97[2] <= stage6_col97[3];
                    stage7_col98[0] <= fa_s6_c97_n57_c;
                    stage7_col98[1] <= fa_s6_c98_n58_s;
                    stage7_col98[2] <= stage6_col98[3];
                    stage7_col99[0] <= fa_s6_c98_n58_c;
                    stage7_col99[1] <= fa_s6_c99_n59_s;
                    stage7_col99[2] <= stage6_col99[3];
                    stage7_col100[0] <= fa_s6_c99_n59_c;
                    stage7_col100[1] <= fa_s6_c100_n60_s;
                    stage7_col100[2] <= stage6_col100[3];
                    stage7_col101[0] <= fa_s6_c100_n60_c;
                    stage7_col101[1] <= fa_s6_c101_n61_s;
                    stage7_col101[2] <= stage6_col101[3];
                    stage7_col102[0] <= fa_s6_c101_n61_c;
                    stage7_col102[1] <= fa_s6_c102_n62_s;
                    stage7_col102[2] <= stage6_col102[3];
                    stage7_col103[0] <= fa_s6_c102_n62_c;
                    stage7_col103[1] <= fa_s6_c103_n63_s;
                    stage7_col103[2] <= stage6_col103[3];
                    stage7_col104[0] <= fa_s6_c103_n63_c;
                    stage7_col104[1] <= fa_s6_c104_n64_s;
                    stage7_col104[2] <= stage6_col104[3];
                    stage7_col105[0] <= fa_s6_c104_n64_c;
                    stage7_col105[1] <= fa_s6_c105_n65_s;
                    stage7_col105[2] <= stage6_col105[3];
                    stage7_col106[0] <= fa_s6_c105_n65_c;
                    stage7_col106[1] <= fa_s6_c106_n66_s;
                    stage7_col106[2] <= stage6_col106[3];
                    stage7_col107[0] <= fa_s6_c106_n66_c;
                    stage7_col107[1] <= fa_s6_c107_n67_s;
                    stage7_col107[2] <= stage6_col107[3];
                    stage7_col108[0] <= fa_s6_c107_n67_c;
                    stage7_col108[1] <= fa_s6_c108_n68_s;
                    stage7_col108[2] <= stage6_col108[3];
                    stage7_col109[0] <= fa_s6_c108_n68_c;
                    stage7_col109[1] <= fa_s6_c109_n69_s;
                    stage7_col109[2] <= stage6_col109[3];
                    stage7_col110[0] <= fa_s6_c109_n69_c;
                    stage7_col110[1] <= fa_s6_c110_n70_s;
                    stage7_col110[2] <= stage6_col110[3];
                    stage7_col111[0] <= fa_s6_c110_n70_c;
                    stage7_col111[1] <= fa_s6_c111_n71_s;
                    stage7_col111[2] <= stage6_col111[3];
                    stage7_col112[0] <= fa_s6_c111_n71_c;
                    stage7_col112[1] <= fa_s6_c112_n72_s;
                    stage7_col112[2] <= stage6_col112[3];
                    stage7_col113[0] <= fa_s6_c112_n72_c;
                    stage7_col113[1] <= fa_s6_c113_n73_s;
                    stage7_col113[2] <= stage6_col113[3];
                    stage7_col114[0] <= fa_s6_c113_n73_c;
                    stage7_col114[1] <= fa_s6_c114_n74_s;
                    stage7_col114[2] <= stage6_col114[3];
                    stage7_col115[0] <= fa_s6_c114_n74_c;
                    stage7_col115[1] <= fa_s6_c115_n75_s;
                    stage7_col115[2] <= stage6_col115[3];
                    stage7_col116[0] <= fa_s6_c115_n75_c;
                    stage7_col116[1] <= fa_s6_c116_n76_s;
                    stage7_col116[2] <= stage6_col116[3];
                    stage7_col117[0] <= fa_s6_c116_n76_c;
                    stage7_col117[1] <= fa_s6_c117_n77_s;
                    stage7_col117[2] <= stage6_col117[3];
                    stage7_col118[0] <= fa_s6_c117_n77_c;
                    stage7_col118[1] <= fa_s6_c118_n78_s;
                    stage7_col118[2] <= stage6_col118[3];
                    stage7_col119[0] <= fa_s6_c118_n78_c;
                    stage7_col119[1] <= fa_s6_c119_n79_s;
                    stage7_col119[2] <= stage6_col119[3];
                    stage7_col120[0] <= fa_s6_c119_n79_c;
                    stage7_col120[1] <= fa_s6_c120_n80_s;
                    stage7_col120[2] <= stage6_col120[3];
                    stage7_col121[0] <= fa_s6_c120_n80_c;
                    stage7_col121[1] <= fa_s6_c121_n81_s;
                    stage7_col121[2] <= stage6_col121[3];
                    stage7_col122[0] <= fa_s6_c121_n81_c;
                    stage7_col122[1] <= fa_s6_c122_n82_s;
                    stage7_col122[2] <= stage6_col122[3];
                    stage7_col123[0] <= fa_s6_c122_n82_c;
                    stage7_col123[1] <= fa_s6_c123_n83_s;
                    stage7_col123[2] <= stage6_col123[3];
                    stage7_col124[0] <= fa_s6_c123_n83_c;
                    stage7_col124[1] <= fa_s6_c124_n84_s;
                    stage7_col124[2] <= stage6_col124[3];
                    stage7_col125[0] <= fa_s6_c124_n84_c;
                    stage7_col125[1] <= fa_s6_c125_n85_s;
                    stage7_col125[2] <= stage6_col125[3];
                    stage7_col126[0] <= fa_s6_c125_n85_c;
                    stage7_col126[1] <= fa_s6_c126_n86_s;
                    stage7_col126[2] <= stage6_col126[3];
                    stage7_col127[0] <= fa_s6_c126_n86_c;
                    stage7_col127[1] <= stage6_col127[0];
                    stage7_col127[2] <= stage6_col127[1];
                    stage7_col127[3] <= stage6_col127[2];
                    stage7_col127[4] <= stage6_col127[3];
                    stage7_col127[5] <= stage6_col127[4];
                    stage7_col127[6] <= stage6_col127[5];
                    stage7_col127[7] <= stage6_col127[6];
                    stage7_col127[8] <= stage6_col127[7];
                    stage7_col127[9] <= stage6_col127[8];
                    stage7_col127[10] <= stage6_col127[9];
                    stage7_col127[11] <= stage6_col127[10];
                    stage7_col127[12] <= stage6_col127[11];
                    stage7_col127[13] <= stage6_col127[12];
                    stage7_col127[14] <= stage6_col127[13];
                    stage7_col127[15] <= stage6_col127[14];
                    stage7_col127[16] <= stage6_col127[15];
                    stage7_col127[17] <= stage6_col127[16];
                    stage7_col127[18] <= stage6_col127[17];
                    stage7_col127[19] <= stage6_col127[18];
                    stage7_col127[20] <= stage6_col127[19];
                    stage7_col127[21] <= stage6_col127[20];
                    stage7_col127[22] <= stage6_col127[21];
                    stage7_col127[23] <= stage6_col127[22];
                    stage7_col127[24] <= stage6_col127[23];
                    stage7_col127[25] <= stage6_col127[24];
                    stage7_col127[26] <= stage6_col127[25];
                    stage7_col127[27] <= stage6_col127[26];
                    stage7_col127[28] <= stage6_col127[27];
                    stage7_col127[29] <= stage6_col127[28];
                    stage7_col127[30] <= stage6_col127[29];
                    stage7_col127[31] <= stage6_col127[29];
                    stage7_col127[32] <= stage6_col127[29];
                    stage7_col127[33] <= stage6_col127[29];
                    stage7_col127[34] <= stage6_col127[29];
                    stage7_col127[35] <= stage6_col127[29];
                    stage7_col127[36] <= stage6_col127[29];
                    stage7_col127[37] <= stage6_col127[29];
                    stage7_col127[38] <= stage6_col127[29];
                    stage7_col127[39] <= stage6_col127[29];
                    stage7_col127[40] <= stage6_col127[29];
                    stage7_col127[41] <= stage6_col127[29];
                    stage7_col127[42] <= stage6_col127[29];
                    stage7_col127[43] <= stage6_col127[29];
                    stage7_col127[44] <= stage6_col127[29];
                    stage7_col127[45] <= stage6_col127[29];
                    stage7_col127[46] <= stage6_col127[29];
                    stage7_col127[47] <= stage6_col127[29];
                    stage7_col127[48] <= stage6_col127[29];
                    stage7_col127[49] <= stage6_col127[29];
                    stage7_col127[50] <= stage6_col127[29];
                    stage7_col127[51] <= stage6_col127[29];
                    stage7_col127[52] <= stage6_col127[29];
                    stage7_col127[53] <= stage6_col127[29];
                    stage7_col127[54] <= stage6_col127[29];
                    stage7_col127[55] <= stage6_col127[29];
                    stage7_col127[56] <= stage6_col127[29];
                    stage7_col127[57] <= stage6_col127[29];
                    stage7_col127[58] <= stage6_col127[29];
                    stage7_col127[59] <= stage6_col127[29];
                    stage7_col127[60] <= stage6_col127[29];
                    stage7_col127[61] <= stage6_col127[29];
                end
            end
        end else begin : gen_stage7_no_pipe
            // Combinational assignment
            always_comb begin
                stage7_col0[0] = stage6_col0[0];
                stage7_col1[0] = stage6_col1[0];
                stage7_col2[0] = stage6_col2[0];
                stage7_col3[0] = stage6_col3[0];
                stage7_col4[0] = stage6_col4[0];
                stage7_col5[0] = stage6_col5[0];
                stage7_col6[0] = ha_s6_c6_n0_s;
                stage7_col7[0] = ha_s6_c6_n0_c;
                stage7_col7[1] = stage6_col7[0];
                stage7_col8[0] = fa_s6_c8_n0_s;
                stage7_col9[0] = fa_s6_c8_n0_c;
                stage7_col9[1] = stage6_col9[0];
                stage7_col9[2] = stage6_col9[1];
                stage7_col10[0] = stage6_col10[0];
                stage7_col10[1] = stage6_col10[1];
                stage7_col11[0] = stage6_col11[0];
                stage7_col11[1] = stage6_col11[1];
                stage7_col12[0] = stage6_col12[0];
                stage7_col12[1] = stage6_col12[1];
                stage7_col13[0] = stage6_col13[0];
                stage7_col13[1] = stage6_col13[1];
                stage7_col14[0] = stage6_col14[0];
                stage7_col14[1] = stage6_col14[1];
                stage7_col15[0] = stage6_col15[0];
                stage7_col15[1] = stage6_col15[1];
                stage7_col16[0] = stage6_col16[0];
                stage7_col16[1] = stage6_col16[1];
                stage7_col17[0] = stage6_col17[0];
                stage7_col17[1] = stage6_col17[1];
                stage7_col18[0] = stage6_col18[0];
                stage7_col18[1] = stage6_col18[1];
                stage7_col19[0] = stage6_col19[0];
                stage7_col19[1] = stage6_col19[1];
                stage7_col20[0] = stage6_col20[0];
                stage7_col20[1] = stage6_col20[1];
                stage7_col21[0] = stage6_col21[0];
                stage7_col21[1] = stage6_col21[1];
                stage7_col22[0] = stage6_col22[0];
                stage7_col22[1] = stage6_col22[1];
                stage7_col23[0] = stage6_col23[0];
                stage7_col23[1] = stage6_col23[1];
                stage7_col24[0] = stage6_col24[0];
                stage7_col24[1] = stage6_col24[1];
                stage7_col25[0] = stage6_col25[0];
                stage7_col25[1] = stage6_col25[1];
                stage7_col26[0] = stage6_col26[0];
                stage7_col26[1] = stage6_col26[1];
                stage7_col27[0] = stage6_col27[0];
                stage7_col27[1] = stage6_col27[1];
                stage7_col28[0] = stage6_col28[0];
                stage7_col28[1] = stage6_col28[1];
                stage7_col29[0] = stage6_col29[0];
                stage7_col29[1] = stage6_col29[1];
                stage7_col30[0] = stage6_col30[0];
                stage7_col30[1] = stage6_col30[1];
                stage7_col31[0] = stage6_col31[0];
                stage7_col31[1] = stage6_col31[1];
                stage7_col32[0] = stage6_col32[0];
                stage7_col32[1] = stage6_col32[1];
                stage7_col33[0] = stage6_col33[0];
                stage7_col33[1] = stage6_col33[1];
                stage7_col34[0] = stage6_col34[0];
                stage7_col34[1] = stage6_col34[1];
                stage7_col35[0] = stage6_col35[0];
                stage7_col35[1] = stage6_col35[1];
                stage7_col36[0] = stage6_col36[0];
                stage7_col36[1] = stage6_col36[1];
                stage7_col37[0] = stage6_col37[0];
                stage7_col37[1] = stage6_col37[1];
                stage7_col38[0] = stage6_col38[0];
                stage7_col38[1] = stage6_col38[1];
                stage7_col39[0] = stage6_col39[0];
                stage7_col39[1] = stage6_col39[1];
                stage7_col40[0] = stage6_col40[0];
                stage7_col40[1] = stage6_col40[1];
                stage7_col41[0] = fa_s6_c41_n1_s;
                stage7_col41[1] = stage6_col41[3];
                stage7_col42[0] = fa_s6_c41_n1_c;
                stage7_col42[1] = fa_s6_c42_n2_s;
                stage7_col43[0] = fa_s6_c42_n2_c;
                stage7_col43[1] = fa_s6_c43_n3_s;
                stage7_col44[0] = fa_s6_c43_n3_c;
                stage7_col44[1] = fa_s6_c44_n4_s;
                stage7_col45[0] = fa_s6_c44_n4_c;
                stage7_col45[1] = fa_s6_c45_n5_s;
                stage7_col46[0] = fa_s6_c45_n5_c;
                stage7_col46[1] = fa_s6_c46_n6_s;
                stage7_col47[0] = fa_s6_c46_n6_c;
                stage7_col47[1] = fa_s6_c47_n7_s;
                stage7_col48[0] = fa_s6_c47_n7_c;
                stage7_col48[1] = fa_s6_c48_n8_s;
                stage7_col49[0] = fa_s6_c48_n8_c;
                stage7_col49[1] = fa_s6_c49_n9_s;
                stage7_col50[0] = fa_s6_c49_n9_c;
                stage7_col50[1] = fa_s6_c50_n10_s;
                stage7_col51[0] = fa_s6_c50_n10_c;
                stage7_col51[1] = fa_s6_c51_n11_s;
                stage7_col52[0] = fa_s6_c51_n11_c;
                stage7_col52[1] = fa_s6_c52_n12_s;
                stage7_col53[0] = fa_s6_c52_n12_c;
                stage7_col53[1] = fa_s6_c53_n13_s;
                stage7_col54[0] = fa_s6_c53_n13_c;
                stage7_col54[1] = fa_s6_c54_n14_s;
                stage7_col55[0] = fa_s6_c54_n14_c;
                stage7_col55[1] = fa_s6_c55_n15_s;
                stage7_col56[0] = fa_s6_c55_n15_c;
                stage7_col56[1] = fa_s6_c56_n16_s;
                stage7_col57[0] = fa_s6_c56_n16_c;
                stage7_col57[1] = fa_s6_c57_n17_s;
                stage7_col58[0] = fa_s6_c57_n17_c;
                stage7_col58[1] = fa_s6_c58_n18_s;
                stage7_col59[0] = fa_s6_c58_n18_c;
                stage7_col59[1] = fa_s6_c59_n19_s;
                stage7_col60[0] = fa_s6_c59_n19_c;
                stage7_col60[1] = fa_s6_c60_n20_s;
                stage7_col60[2] = stage6_col60[3];
                stage7_col61[0] = fa_s6_c60_n20_c;
                stage7_col61[1] = fa_s6_c61_n21_s;
                stage7_col61[2] = stage6_col61[3];
                stage7_col62[0] = fa_s6_c61_n21_c;
                stage7_col62[1] = fa_s6_c62_n22_s;
                stage7_col62[2] = stage6_col62[3];
                stage7_col63[0] = fa_s6_c62_n22_c;
                stage7_col63[1] = fa_s6_c63_n23_s;
                stage7_col63[2] = stage6_col63[3];
                stage7_col64[0] = fa_s6_c63_n23_c;
                stage7_col64[1] = fa_s6_c64_n24_s;
                stage7_col64[2] = stage6_col64[3];
                stage7_col65[0] = fa_s6_c64_n24_c;
                stage7_col65[1] = fa_s6_c65_n25_s;
                stage7_col65[2] = stage6_col65[3];
                stage7_col66[0] = fa_s6_c65_n25_c;
                stage7_col66[1] = fa_s6_c66_n26_s;
                stage7_col66[2] = stage6_col66[3];
                stage7_col67[0] = fa_s6_c66_n26_c;
                stage7_col67[1] = fa_s6_c67_n27_s;
                stage7_col67[2] = stage6_col67[3];
                stage7_col68[0] = fa_s6_c67_n27_c;
                stage7_col68[1] = fa_s6_c68_n28_s;
                stage7_col68[2] = stage6_col68[3];
                stage7_col69[0] = fa_s6_c68_n28_c;
                stage7_col69[1] = fa_s6_c69_n29_s;
                stage7_col69[2] = stage6_col69[3];
                stage7_col70[0] = fa_s6_c69_n29_c;
                stage7_col70[1] = fa_s6_c70_n30_s;
                stage7_col70[2] = stage6_col70[3];
                stage7_col71[0] = fa_s6_c70_n30_c;
                stage7_col71[1] = fa_s6_c71_n31_s;
                stage7_col71[2] = stage6_col71[3];
                stage7_col72[0] = fa_s6_c71_n31_c;
                stage7_col72[1] = fa_s6_c72_n32_s;
                stage7_col72[2] = stage6_col72[3];
                stage7_col73[0] = fa_s6_c72_n32_c;
                stage7_col73[1] = fa_s6_c73_n33_s;
                stage7_col73[2] = stage6_col73[3];
                stage7_col74[0] = fa_s6_c73_n33_c;
                stage7_col74[1] = fa_s6_c74_n34_s;
                stage7_col74[2] = stage6_col74[3];
                stage7_col75[0] = fa_s6_c74_n34_c;
                stage7_col75[1] = fa_s6_c75_n35_s;
                stage7_col75[2] = stage6_col75[3];
                stage7_col76[0] = fa_s6_c75_n35_c;
                stage7_col76[1] = fa_s6_c76_n36_s;
                stage7_col76[2] = stage6_col76[3];
                stage7_col77[0] = fa_s6_c76_n36_c;
                stage7_col77[1] = fa_s6_c77_n37_s;
                stage7_col77[2] = stage6_col77[3];
                stage7_col78[0] = fa_s6_c77_n37_c;
                stage7_col78[1] = fa_s6_c78_n38_s;
                stage7_col78[2] = stage6_col78[3];
                stage7_col79[0] = fa_s6_c78_n38_c;
                stage7_col79[1] = fa_s6_c79_n39_s;
                stage7_col79[2] = stage6_col79[3];
                stage7_col80[0] = fa_s6_c79_n39_c;
                stage7_col80[1] = fa_s6_c80_n40_s;
                stage7_col80[2] = stage6_col80[3];
                stage7_col81[0] = fa_s6_c80_n40_c;
                stage7_col81[1] = fa_s6_c81_n41_s;
                stage7_col81[2] = stage6_col81[3];
                stage7_col82[0] = fa_s6_c81_n41_c;
                stage7_col82[1] = fa_s6_c82_n42_s;
                stage7_col82[2] = stage6_col82[3];
                stage7_col83[0] = fa_s6_c82_n42_c;
                stage7_col83[1] = fa_s6_c83_n43_s;
                stage7_col83[2] = stage6_col83[3];
                stage7_col84[0] = fa_s6_c83_n43_c;
                stage7_col84[1] = fa_s6_c84_n44_s;
                stage7_col84[2] = stage6_col84[3];
                stage7_col85[0] = fa_s6_c84_n44_c;
                stage7_col85[1] = fa_s6_c85_n45_s;
                stage7_col85[2] = stage6_col85[3];
                stage7_col86[0] = fa_s6_c85_n45_c;
                stage7_col86[1] = fa_s6_c86_n46_s;
                stage7_col86[2] = stage6_col86[3];
                stage7_col87[0] = fa_s6_c86_n46_c;
                stage7_col87[1] = fa_s6_c87_n47_s;
                stage7_col87[2] = stage6_col87[3];
                stage7_col88[0] = fa_s6_c87_n47_c;
                stage7_col88[1] = fa_s6_c88_n48_s;
                stage7_col88[2] = stage6_col88[3];
                stage7_col89[0] = fa_s6_c88_n48_c;
                stage7_col89[1] = fa_s6_c89_n49_s;
                stage7_col89[2] = stage6_col89[3];
                stage7_col90[0] = fa_s6_c89_n49_c;
                stage7_col90[1] = fa_s6_c90_n50_s;
                stage7_col90[2] = stage6_col90[3];
                stage7_col91[0] = fa_s6_c90_n50_c;
                stage7_col91[1] = fa_s6_c91_n51_s;
                stage7_col91[2] = stage6_col91[3];
                stage7_col92[0] = fa_s6_c91_n51_c;
                stage7_col92[1] = fa_s6_c92_n52_s;
                stage7_col92[2] = stage6_col92[3];
                stage7_col93[0] = fa_s6_c92_n52_c;
                stage7_col93[1] = fa_s6_c93_n53_s;
                stage7_col93[2] = stage6_col93[3];
                stage7_col94[0] = fa_s6_c93_n53_c;
                stage7_col94[1] = fa_s6_c94_n54_s;
                stage7_col94[2] = stage6_col94[3];
                stage7_col95[0] = fa_s6_c94_n54_c;
                stage7_col95[1] = fa_s6_c95_n55_s;
                stage7_col95[2] = stage6_col95[3];
                stage7_col96[0] = fa_s6_c95_n55_c;
                stage7_col96[1] = fa_s6_c96_n56_s;
                stage7_col96[2] = stage6_col96[3];
                stage7_col97[0] = fa_s6_c96_n56_c;
                stage7_col97[1] = fa_s6_c97_n57_s;
                stage7_col97[2] = stage6_col97[3];
                stage7_col98[0] = fa_s6_c97_n57_c;
                stage7_col98[1] = fa_s6_c98_n58_s;
                stage7_col98[2] = stage6_col98[3];
                stage7_col99[0] = fa_s6_c98_n58_c;
                stage7_col99[1] = fa_s6_c99_n59_s;
                stage7_col99[2] = stage6_col99[3];
                stage7_col100[0] = fa_s6_c99_n59_c;
                stage7_col100[1] = fa_s6_c100_n60_s;
                stage7_col100[2] = stage6_col100[3];
                stage7_col101[0] = fa_s6_c100_n60_c;
                stage7_col101[1] = fa_s6_c101_n61_s;
                stage7_col101[2] = stage6_col101[3];
                stage7_col102[0] = fa_s6_c101_n61_c;
                stage7_col102[1] = fa_s6_c102_n62_s;
                stage7_col102[2] = stage6_col102[3];
                stage7_col103[0] = fa_s6_c102_n62_c;
                stage7_col103[1] = fa_s6_c103_n63_s;
                stage7_col103[2] = stage6_col103[3];
                stage7_col104[0] = fa_s6_c103_n63_c;
                stage7_col104[1] = fa_s6_c104_n64_s;
                stage7_col104[2] = stage6_col104[3];
                stage7_col105[0] = fa_s6_c104_n64_c;
                stage7_col105[1] = fa_s6_c105_n65_s;
                stage7_col105[2] = stage6_col105[3];
                stage7_col106[0] = fa_s6_c105_n65_c;
                stage7_col106[1] = fa_s6_c106_n66_s;
                stage7_col106[2] = stage6_col106[3];
                stage7_col107[0] = fa_s6_c106_n66_c;
                stage7_col107[1] = fa_s6_c107_n67_s;
                stage7_col107[2] = stage6_col107[3];
                stage7_col108[0] = fa_s6_c107_n67_c;
                stage7_col108[1] = fa_s6_c108_n68_s;
                stage7_col108[2] = stage6_col108[3];
                stage7_col109[0] = fa_s6_c108_n68_c;
                stage7_col109[1] = fa_s6_c109_n69_s;
                stage7_col109[2] = stage6_col109[3];
                stage7_col110[0] = fa_s6_c109_n69_c;
                stage7_col110[1] = fa_s6_c110_n70_s;
                stage7_col110[2] = stage6_col110[3];
                stage7_col111[0] = fa_s6_c110_n70_c;
                stage7_col111[1] = fa_s6_c111_n71_s;
                stage7_col111[2] = stage6_col111[3];
                stage7_col112[0] = fa_s6_c111_n71_c;
                stage7_col112[1] = fa_s6_c112_n72_s;
                stage7_col112[2] = stage6_col112[3];
                stage7_col113[0] = fa_s6_c112_n72_c;
                stage7_col113[1] = fa_s6_c113_n73_s;
                stage7_col113[2] = stage6_col113[3];
                stage7_col114[0] = fa_s6_c113_n73_c;
                stage7_col114[1] = fa_s6_c114_n74_s;
                stage7_col114[2] = stage6_col114[3];
                stage7_col115[0] = fa_s6_c114_n74_c;
                stage7_col115[1] = fa_s6_c115_n75_s;
                stage7_col115[2] = stage6_col115[3];
                stage7_col116[0] = fa_s6_c115_n75_c;
                stage7_col116[1] = fa_s6_c116_n76_s;
                stage7_col116[2] = stage6_col116[3];
                stage7_col117[0] = fa_s6_c116_n76_c;
                stage7_col117[1] = fa_s6_c117_n77_s;
                stage7_col117[2] = stage6_col117[3];
                stage7_col118[0] = fa_s6_c117_n77_c;
                stage7_col118[1] = fa_s6_c118_n78_s;
                stage7_col118[2] = stage6_col118[3];
                stage7_col119[0] = fa_s6_c118_n78_c;
                stage7_col119[1] = fa_s6_c119_n79_s;
                stage7_col119[2] = stage6_col119[3];
                stage7_col120[0] = fa_s6_c119_n79_c;
                stage7_col120[1] = fa_s6_c120_n80_s;
                stage7_col120[2] = stage6_col120[3];
                stage7_col121[0] = fa_s6_c120_n80_c;
                stage7_col121[1] = fa_s6_c121_n81_s;
                stage7_col121[2] = stage6_col121[3];
                stage7_col122[0] = fa_s6_c121_n81_c;
                stage7_col122[1] = fa_s6_c122_n82_s;
                stage7_col122[2] = stage6_col122[3];
                stage7_col123[0] = fa_s6_c122_n82_c;
                stage7_col123[1] = fa_s6_c123_n83_s;
                stage7_col123[2] = stage6_col123[3];
                stage7_col124[0] = fa_s6_c123_n83_c;
                stage7_col124[1] = fa_s6_c124_n84_s;
                stage7_col124[2] = stage6_col124[3];
                stage7_col125[0] = fa_s6_c124_n84_c;
                stage7_col125[1] = fa_s6_c125_n85_s;
                stage7_col125[2] = stage6_col125[3];
                stage7_col126[0] = fa_s6_c125_n85_c;
                stage7_col126[1] = fa_s6_c126_n86_s;
                stage7_col126[2] = stage6_col126[3];
                stage7_col127[0] = fa_s6_c126_n86_c;
                stage7_col127[1] = stage6_col127[0];
                stage7_col127[2] = stage6_col127[1];
                stage7_col127[3] = stage6_col127[2];
                stage7_col127[4] = stage6_col127[3];
                stage7_col127[5] = stage6_col127[4];
                stage7_col127[6] = stage6_col127[5];
                stage7_col127[7] = stage6_col127[6];
                stage7_col127[8] = stage6_col127[7];
                stage7_col127[9] = stage6_col127[8];
                stage7_col127[10] = stage6_col127[9];
                stage7_col127[11] = stage6_col127[10];
                stage7_col127[12] = stage6_col127[11];
                stage7_col127[13] = stage6_col127[12];
                stage7_col127[14] = stage6_col127[13];
                stage7_col127[15] = stage6_col127[14];
                stage7_col127[16] = stage6_col127[15];
                stage7_col127[17] = stage6_col127[16];
                stage7_col127[18] = stage6_col127[17];
                stage7_col127[19] = stage6_col127[18];
                stage7_col127[20] = stage6_col127[19];
                stage7_col127[21] = stage6_col127[20];
                stage7_col127[22] = stage6_col127[21];
                stage7_col127[23] = stage6_col127[22];
                stage7_col127[24] = stage6_col127[23];
                stage7_col127[25] = stage6_col127[24];
                stage7_col127[26] = stage6_col127[25];
                stage7_col127[27] = stage6_col127[26];
                stage7_col127[28] = stage6_col127[27];
                stage7_col127[29] = stage6_col127[28];
                stage7_col127[30] = stage6_col127[29];
                stage7_col127[31] = stage6_col127[29];
                stage7_col127[32] = stage6_col127[29];
                stage7_col127[33] = stage6_col127[29];
                stage7_col127[34] = stage6_col127[29];
                stage7_col127[35] = stage6_col127[29];
                stage7_col127[36] = stage6_col127[29];
                stage7_col127[37] = stage6_col127[29];
                stage7_col127[38] = stage6_col127[29];
                stage7_col127[39] = stage6_col127[29];
                stage7_col127[40] = stage6_col127[29];
                stage7_col127[41] = stage6_col127[29];
                stage7_col127[42] = stage6_col127[29];
                stage7_col127[43] = stage6_col127[29];
                stage7_col127[44] = stage6_col127[29];
                stage7_col127[45] = stage6_col127[29];
                stage7_col127[46] = stage6_col127[29];
                stage7_col127[47] = stage6_col127[29];
                stage7_col127[48] = stage6_col127[29];
                stage7_col127[49] = stage6_col127[29];
                stage7_col127[50] = stage6_col127[29];
                stage7_col127[51] = stage6_col127[29];
                stage7_col127[52] = stage6_col127[29];
                stage7_col127[53] = stage6_col127[29];
                stage7_col127[54] = stage6_col127[29];
                stage7_col127[55] = stage6_col127[29];
                stage7_col127[56] = stage6_col127[29];
                stage7_col127[57] = stage6_col127[29];
                stage7_col127[58] = stage6_col127[29];
                stage7_col127[59] = stage6_col127[29];
                stage7_col127[60] = stage6_col127[29];
                stage7_col127[61] = stage6_col127[29];
            end
        end
    endgenerate

    // Stage 8: Reduction
    fa fa_s7_c9_n0 (
        .a(stage7_col9[0]),
        .b(stage7_col9[1]),
        .c_in(stage7_col9[2]),
        .s(fa_s7_c9_n0_s),
        .c_out(fa_s7_c9_n0_c)
    );

    fa fa_s7_c60_n1 (
        .a(stage7_col60[0]),
        .b(stage7_col60[1]),
        .c_in(stage7_col60[2]),
        .s(fa_s7_c60_n1_s),
        .c_out(fa_s7_c60_n1_c)
    );

    fa fa_s7_c61_n2 (
        .a(stage7_col61[0]),
        .b(stage7_col61[1]),
        .c_in(stage7_col61[2]),
        .s(fa_s7_c61_n2_s),
        .c_out(fa_s7_c61_n2_c)
    );

    fa fa_s7_c62_n3 (
        .a(stage7_col62[0]),
        .b(stage7_col62[1]),
        .c_in(stage7_col62[2]),
        .s(fa_s7_c62_n3_s),
        .c_out(fa_s7_c62_n3_c)
    );

    fa fa_s7_c63_n4 (
        .a(stage7_col63[0]),
        .b(stage7_col63[1]),
        .c_in(stage7_col63[2]),
        .s(fa_s7_c63_n4_s),
        .c_out(fa_s7_c63_n4_c)
    );

    fa fa_s7_c64_n5 (
        .a(stage7_col64[0]),
        .b(stage7_col64[1]),
        .c_in(stage7_col64[2]),
        .s(fa_s7_c64_n5_s),
        .c_out(fa_s7_c64_n5_c)
    );

    fa fa_s7_c65_n6 (
        .a(stage7_col65[0]),
        .b(stage7_col65[1]),
        .c_in(stage7_col65[2]),
        .s(fa_s7_c65_n6_s),
        .c_out(fa_s7_c65_n6_c)
    );

    fa fa_s7_c66_n7 (
        .a(stage7_col66[0]),
        .b(stage7_col66[1]),
        .c_in(stage7_col66[2]),
        .s(fa_s7_c66_n7_s),
        .c_out(fa_s7_c66_n7_c)
    );

    fa fa_s7_c67_n8 (
        .a(stage7_col67[0]),
        .b(stage7_col67[1]),
        .c_in(stage7_col67[2]),
        .s(fa_s7_c67_n8_s),
        .c_out(fa_s7_c67_n8_c)
    );

    fa fa_s7_c68_n9 (
        .a(stage7_col68[0]),
        .b(stage7_col68[1]),
        .c_in(stage7_col68[2]),
        .s(fa_s7_c68_n9_s),
        .c_out(fa_s7_c68_n9_c)
    );

    fa fa_s7_c69_n10 (
        .a(stage7_col69[0]),
        .b(stage7_col69[1]),
        .c_in(stage7_col69[2]),
        .s(fa_s7_c69_n10_s),
        .c_out(fa_s7_c69_n10_c)
    );

    fa fa_s7_c70_n11 (
        .a(stage7_col70[0]),
        .b(stage7_col70[1]),
        .c_in(stage7_col70[2]),
        .s(fa_s7_c70_n11_s),
        .c_out(fa_s7_c70_n11_c)
    );

    fa fa_s7_c71_n12 (
        .a(stage7_col71[0]),
        .b(stage7_col71[1]),
        .c_in(stage7_col71[2]),
        .s(fa_s7_c71_n12_s),
        .c_out(fa_s7_c71_n12_c)
    );

    fa fa_s7_c72_n13 (
        .a(stage7_col72[0]),
        .b(stage7_col72[1]),
        .c_in(stage7_col72[2]),
        .s(fa_s7_c72_n13_s),
        .c_out(fa_s7_c72_n13_c)
    );

    fa fa_s7_c73_n14 (
        .a(stage7_col73[0]),
        .b(stage7_col73[1]),
        .c_in(stage7_col73[2]),
        .s(fa_s7_c73_n14_s),
        .c_out(fa_s7_c73_n14_c)
    );

    fa fa_s7_c74_n15 (
        .a(stage7_col74[0]),
        .b(stage7_col74[1]),
        .c_in(stage7_col74[2]),
        .s(fa_s7_c74_n15_s),
        .c_out(fa_s7_c74_n15_c)
    );

    fa fa_s7_c75_n16 (
        .a(stage7_col75[0]),
        .b(stage7_col75[1]),
        .c_in(stage7_col75[2]),
        .s(fa_s7_c75_n16_s),
        .c_out(fa_s7_c75_n16_c)
    );

    fa fa_s7_c76_n17 (
        .a(stage7_col76[0]),
        .b(stage7_col76[1]),
        .c_in(stage7_col76[2]),
        .s(fa_s7_c76_n17_s),
        .c_out(fa_s7_c76_n17_c)
    );

    fa fa_s7_c77_n18 (
        .a(stage7_col77[0]),
        .b(stage7_col77[1]),
        .c_in(stage7_col77[2]),
        .s(fa_s7_c77_n18_s),
        .c_out(fa_s7_c77_n18_c)
    );

    fa fa_s7_c78_n19 (
        .a(stage7_col78[0]),
        .b(stage7_col78[1]),
        .c_in(stage7_col78[2]),
        .s(fa_s7_c78_n19_s),
        .c_out(fa_s7_c78_n19_c)
    );

    fa fa_s7_c79_n20 (
        .a(stage7_col79[0]),
        .b(stage7_col79[1]),
        .c_in(stage7_col79[2]),
        .s(fa_s7_c79_n20_s),
        .c_out(fa_s7_c79_n20_c)
    );

    fa fa_s7_c80_n21 (
        .a(stage7_col80[0]),
        .b(stage7_col80[1]),
        .c_in(stage7_col80[2]),
        .s(fa_s7_c80_n21_s),
        .c_out(fa_s7_c80_n21_c)
    );

    fa fa_s7_c81_n22 (
        .a(stage7_col81[0]),
        .b(stage7_col81[1]),
        .c_in(stage7_col81[2]),
        .s(fa_s7_c81_n22_s),
        .c_out(fa_s7_c81_n22_c)
    );

    fa fa_s7_c82_n23 (
        .a(stage7_col82[0]),
        .b(stage7_col82[1]),
        .c_in(stage7_col82[2]),
        .s(fa_s7_c82_n23_s),
        .c_out(fa_s7_c82_n23_c)
    );

    fa fa_s7_c83_n24 (
        .a(stage7_col83[0]),
        .b(stage7_col83[1]),
        .c_in(stage7_col83[2]),
        .s(fa_s7_c83_n24_s),
        .c_out(fa_s7_c83_n24_c)
    );

    fa fa_s7_c84_n25 (
        .a(stage7_col84[0]),
        .b(stage7_col84[1]),
        .c_in(stage7_col84[2]),
        .s(fa_s7_c84_n25_s),
        .c_out(fa_s7_c84_n25_c)
    );

    fa fa_s7_c85_n26 (
        .a(stage7_col85[0]),
        .b(stage7_col85[1]),
        .c_in(stage7_col85[2]),
        .s(fa_s7_c85_n26_s),
        .c_out(fa_s7_c85_n26_c)
    );

    fa fa_s7_c86_n27 (
        .a(stage7_col86[0]),
        .b(stage7_col86[1]),
        .c_in(stage7_col86[2]),
        .s(fa_s7_c86_n27_s),
        .c_out(fa_s7_c86_n27_c)
    );

    fa fa_s7_c87_n28 (
        .a(stage7_col87[0]),
        .b(stage7_col87[1]),
        .c_in(stage7_col87[2]),
        .s(fa_s7_c87_n28_s),
        .c_out(fa_s7_c87_n28_c)
    );

    fa fa_s7_c88_n29 (
        .a(stage7_col88[0]),
        .b(stage7_col88[1]),
        .c_in(stage7_col88[2]),
        .s(fa_s7_c88_n29_s),
        .c_out(fa_s7_c88_n29_c)
    );

    fa fa_s7_c89_n30 (
        .a(stage7_col89[0]),
        .b(stage7_col89[1]),
        .c_in(stage7_col89[2]),
        .s(fa_s7_c89_n30_s),
        .c_out(fa_s7_c89_n30_c)
    );

    fa fa_s7_c90_n31 (
        .a(stage7_col90[0]),
        .b(stage7_col90[1]),
        .c_in(stage7_col90[2]),
        .s(fa_s7_c90_n31_s),
        .c_out(fa_s7_c90_n31_c)
    );

    fa fa_s7_c91_n32 (
        .a(stage7_col91[0]),
        .b(stage7_col91[1]),
        .c_in(stage7_col91[2]),
        .s(fa_s7_c91_n32_s),
        .c_out(fa_s7_c91_n32_c)
    );

    fa fa_s7_c92_n33 (
        .a(stage7_col92[0]),
        .b(stage7_col92[1]),
        .c_in(stage7_col92[2]),
        .s(fa_s7_c92_n33_s),
        .c_out(fa_s7_c92_n33_c)
    );

    fa fa_s7_c93_n34 (
        .a(stage7_col93[0]),
        .b(stage7_col93[1]),
        .c_in(stage7_col93[2]),
        .s(fa_s7_c93_n34_s),
        .c_out(fa_s7_c93_n34_c)
    );

    fa fa_s7_c94_n35 (
        .a(stage7_col94[0]),
        .b(stage7_col94[1]),
        .c_in(stage7_col94[2]),
        .s(fa_s7_c94_n35_s),
        .c_out(fa_s7_c94_n35_c)
    );

    fa fa_s7_c95_n36 (
        .a(stage7_col95[0]),
        .b(stage7_col95[1]),
        .c_in(stage7_col95[2]),
        .s(fa_s7_c95_n36_s),
        .c_out(fa_s7_c95_n36_c)
    );

    fa fa_s7_c96_n37 (
        .a(stage7_col96[0]),
        .b(stage7_col96[1]),
        .c_in(stage7_col96[2]),
        .s(fa_s7_c96_n37_s),
        .c_out(fa_s7_c96_n37_c)
    );

    fa fa_s7_c97_n38 (
        .a(stage7_col97[0]),
        .b(stage7_col97[1]),
        .c_in(stage7_col97[2]),
        .s(fa_s7_c97_n38_s),
        .c_out(fa_s7_c97_n38_c)
    );

    fa fa_s7_c98_n39 (
        .a(stage7_col98[0]),
        .b(stage7_col98[1]),
        .c_in(stage7_col98[2]),
        .s(fa_s7_c98_n39_s),
        .c_out(fa_s7_c98_n39_c)
    );

    fa fa_s7_c99_n40 (
        .a(stage7_col99[0]),
        .b(stage7_col99[1]),
        .c_in(stage7_col99[2]),
        .s(fa_s7_c99_n40_s),
        .c_out(fa_s7_c99_n40_c)
    );

    fa fa_s7_c100_n41 (
        .a(stage7_col100[0]),
        .b(stage7_col100[1]),
        .c_in(stage7_col100[2]),
        .s(fa_s7_c100_n41_s),
        .c_out(fa_s7_c100_n41_c)
    );

    fa fa_s7_c101_n42 (
        .a(stage7_col101[0]),
        .b(stage7_col101[1]),
        .c_in(stage7_col101[2]),
        .s(fa_s7_c101_n42_s),
        .c_out(fa_s7_c101_n42_c)
    );

    fa fa_s7_c102_n43 (
        .a(stage7_col102[0]),
        .b(stage7_col102[1]),
        .c_in(stage7_col102[2]),
        .s(fa_s7_c102_n43_s),
        .c_out(fa_s7_c102_n43_c)
    );

    fa fa_s7_c103_n44 (
        .a(stage7_col103[0]),
        .b(stage7_col103[1]),
        .c_in(stage7_col103[2]),
        .s(fa_s7_c103_n44_s),
        .c_out(fa_s7_c103_n44_c)
    );

    fa fa_s7_c104_n45 (
        .a(stage7_col104[0]),
        .b(stage7_col104[1]),
        .c_in(stage7_col104[2]),
        .s(fa_s7_c104_n45_s),
        .c_out(fa_s7_c104_n45_c)
    );

    fa fa_s7_c105_n46 (
        .a(stage7_col105[0]),
        .b(stage7_col105[1]),
        .c_in(stage7_col105[2]),
        .s(fa_s7_c105_n46_s),
        .c_out(fa_s7_c105_n46_c)
    );

    fa fa_s7_c106_n47 (
        .a(stage7_col106[0]),
        .b(stage7_col106[1]),
        .c_in(stage7_col106[2]),
        .s(fa_s7_c106_n47_s),
        .c_out(fa_s7_c106_n47_c)
    );

    fa fa_s7_c107_n48 (
        .a(stage7_col107[0]),
        .b(stage7_col107[1]),
        .c_in(stage7_col107[2]),
        .s(fa_s7_c107_n48_s),
        .c_out(fa_s7_c107_n48_c)
    );

    fa fa_s7_c108_n49 (
        .a(stage7_col108[0]),
        .b(stage7_col108[1]),
        .c_in(stage7_col108[2]),
        .s(fa_s7_c108_n49_s),
        .c_out(fa_s7_c108_n49_c)
    );

    fa fa_s7_c109_n50 (
        .a(stage7_col109[0]),
        .b(stage7_col109[1]),
        .c_in(stage7_col109[2]),
        .s(fa_s7_c109_n50_s),
        .c_out(fa_s7_c109_n50_c)
    );

    fa fa_s7_c110_n51 (
        .a(stage7_col110[0]),
        .b(stage7_col110[1]),
        .c_in(stage7_col110[2]),
        .s(fa_s7_c110_n51_s),
        .c_out(fa_s7_c110_n51_c)
    );

    fa fa_s7_c111_n52 (
        .a(stage7_col111[0]),
        .b(stage7_col111[1]),
        .c_in(stage7_col111[2]),
        .s(fa_s7_c111_n52_s),
        .c_out(fa_s7_c111_n52_c)
    );

    fa fa_s7_c112_n53 (
        .a(stage7_col112[0]),
        .b(stage7_col112[1]),
        .c_in(stage7_col112[2]),
        .s(fa_s7_c112_n53_s),
        .c_out(fa_s7_c112_n53_c)
    );

    fa fa_s7_c113_n54 (
        .a(stage7_col113[0]),
        .b(stage7_col113[1]),
        .c_in(stage7_col113[2]),
        .s(fa_s7_c113_n54_s),
        .c_out(fa_s7_c113_n54_c)
    );

    fa fa_s7_c114_n55 (
        .a(stage7_col114[0]),
        .b(stage7_col114[1]),
        .c_in(stage7_col114[2]),
        .s(fa_s7_c114_n55_s),
        .c_out(fa_s7_c114_n55_c)
    );

    fa fa_s7_c115_n56 (
        .a(stage7_col115[0]),
        .b(stage7_col115[1]),
        .c_in(stage7_col115[2]),
        .s(fa_s7_c115_n56_s),
        .c_out(fa_s7_c115_n56_c)
    );

    fa fa_s7_c116_n57 (
        .a(stage7_col116[0]),
        .b(stage7_col116[1]),
        .c_in(stage7_col116[2]),
        .s(fa_s7_c116_n57_s),
        .c_out(fa_s7_c116_n57_c)
    );

    fa fa_s7_c117_n58 (
        .a(stage7_col117[0]),
        .b(stage7_col117[1]),
        .c_in(stage7_col117[2]),
        .s(fa_s7_c117_n58_s),
        .c_out(fa_s7_c117_n58_c)
    );

    fa fa_s7_c118_n59 (
        .a(stage7_col118[0]),
        .b(stage7_col118[1]),
        .c_in(stage7_col118[2]),
        .s(fa_s7_c118_n59_s),
        .c_out(fa_s7_c118_n59_c)
    );

    fa fa_s7_c119_n60 (
        .a(stage7_col119[0]),
        .b(stage7_col119[1]),
        .c_in(stage7_col119[2]),
        .s(fa_s7_c119_n60_s),
        .c_out(fa_s7_c119_n60_c)
    );

    fa fa_s7_c120_n61 (
        .a(stage7_col120[0]),
        .b(stage7_col120[1]),
        .c_in(stage7_col120[2]),
        .s(fa_s7_c120_n61_s),
        .c_out(fa_s7_c120_n61_c)
    );

    fa fa_s7_c121_n62 (
        .a(stage7_col121[0]),
        .b(stage7_col121[1]),
        .c_in(stage7_col121[2]),
        .s(fa_s7_c121_n62_s),
        .c_out(fa_s7_c121_n62_c)
    );

    fa fa_s7_c122_n63 (
        .a(stage7_col122[0]),
        .b(stage7_col122[1]),
        .c_in(stage7_col122[2]),
        .s(fa_s7_c122_n63_s),
        .c_out(fa_s7_c122_n63_c)
    );

    fa fa_s7_c123_n64 (
        .a(stage7_col123[0]),
        .b(stage7_col123[1]),
        .c_in(stage7_col123[2]),
        .s(fa_s7_c123_n64_s),
        .c_out(fa_s7_c123_n64_c)
    );

    fa fa_s7_c124_n65 (
        .a(stage7_col124[0]),
        .b(stage7_col124[1]),
        .c_in(stage7_col124[2]),
        .s(fa_s7_c124_n65_s),
        .c_out(fa_s7_c124_n65_c)
    );

    fa fa_s7_c125_n66 (
        .a(stage7_col125[0]),
        .b(stage7_col125[1]),
        .c_in(stage7_col125[2]),
        .s(fa_s7_c125_n66_s),
        .c_out(fa_s7_c125_n66_c)
    );

    fa fa_s7_c126_n67 (
        .a(stage7_col126[0]),
        .b(stage7_col126[1]),
        .c_in(stage7_col126[2]),
        .s(fa_s7_c126_n67_s),
        .c_out(fa_s7_c126_n67_c)
    );

    ha ha_s7_c7_n0 (
        .a(stage7_col7[0]),
        .b(stage7_col7[1]),
        .s(ha_s7_c7_n0_s),
        .c_out(ha_s7_c7_n0_c)
    );

    ha ha_s7_c10_n1 (
        .a(stage7_col10[0]),
        .b(stage7_col10[1]),
        .s(ha_s7_c10_n1_s),
        .c_out(ha_s7_c10_n1_c)
    );

    ha ha_s7_c11_n2 (
        .a(stage7_col11[0]),
        .b(stage7_col11[1]),
        .s(ha_s7_c11_n2_s),
        .c_out(ha_s7_c11_n2_c)
    );

    ha ha_s7_c12_n3 (
        .a(stage7_col12[0]),
        .b(stage7_col12[1]),
        .s(ha_s7_c12_n3_s),
        .c_out(ha_s7_c12_n3_c)
    );

    ha ha_s7_c13_n4 (
        .a(stage7_col13[0]),
        .b(stage7_col13[1]),
        .s(ha_s7_c13_n4_s),
        .c_out(ha_s7_c13_n4_c)
    );

    ha ha_s7_c14_n5 (
        .a(stage7_col14[0]),
        .b(stage7_col14[1]),
        .s(ha_s7_c14_n5_s),
        .c_out(ha_s7_c14_n5_c)
    );

    ha ha_s7_c15_n6 (
        .a(stage7_col15[0]),
        .b(stage7_col15[1]),
        .s(ha_s7_c15_n6_s),
        .c_out(ha_s7_c15_n6_c)
    );

    ha ha_s7_c16_n7 (
        .a(stage7_col16[0]),
        .b(stage7_col16[1]),
        .s(ha_s7_c16_n7_s),
        .c_out(ha_s7_c16_n7_c)
    );

    ha ha_s7_c17_n8 (
        .a(stage7_col17[0]),
        .b(stage7_col17[1]),
        .s(ha_s7_c17_n8_s),
        .c_out(ha_s7_c17_n8_c)
    );

    ha ha_s7_c18_n9 (
        .a(stage7_col18[0]),
        .b(stage7_col18[1]),
        .s(ha_s7_c18_n9_s),
        .c_out(ha_s7_c18_n9_c)
    );

    ha ha_s7_c19_n10 (
        .a(stage7_col19[0]),
        .b(stage7_col19[1]),
        .s(ha_s7_c19_n10_s),
        .c_out(ha_s7_c19_n10_c)
    );

    ha ha_s7_c20_n11 (
        .a(stage7_col20[0]),
        .b(stage7_col20[1]),
        .s(ha_s7_c20_n11_s),
        .c_out(ha_s7_c20_n11_c)
    );

    ha ha_s7_c21_n12 (
        .a(stage7_col21[0]),
        .b(stage7_col21[1]),
        .s(ha_s7_c21_n12_s),
        .c_out(ha_s7_c21_n12_c)
    );

    ha ha_s7_c22_n13 (
        .a(stage7_col22[0]),
        .b(stage7_col22[1]),
        .s(ha_s7_c22_n13_s),
        .c_out(ha_s7_c22_n13_c)
    );

    ha ha_s7_c23_n14 (
        .a(stage7_col23[0]),
        .b(stage7_col23[1]),
        .s(ha_s7_c23_n14_s),
        .c_out(ha_s7_c23_n14_c)
    );

    ha ha_s7_c24_n15 (
        .a(stage7_col24[0]),
        .b(stage7_col24[1]),
        .s(ha_s7_c24_n15_s),
        .c_out(ha_s7_c24_n15_c)
    );

    ha ha_s7_c25_n16 (
        .a(stage7_col25[0]),
        .b(stage7_col25[1]),
        .s(ha_s7_c25_n16_s),
        .c_out(ha_s7_c25_n16_c)
    );

    ha ha_s7_c26_n17 (
        .a(stage7_col26[0]),
        .b(stage7_col26[1]),
        .s(ha_s7_c26_n17_s),
        .c_out(ha_s7_c26_n17_c)
    );

    ha ha_s7_c27_n18 (
        .a(stage7_col27[0]),
        .b(stage7_col27[1]),
        .s(ha_s7_c27_n18_s),
        .c_out(ha_s7_c27_n18_c)
    );

    ha ha_s7_c28_n19 (
        .a(stage7_col28[0]),
        .b(stage7_col28[1]),
        .s(ha_s7_c28_n19_s),
        .c_out(ha_s7_c28_n19_c)
    );

    ha ha_s7_c29_n20 (
        .a(stage7_col29[0]),
        .b(stage7_col29[1]),
        .s(ha_s7_c29_n20_s),
        .c_out(ha_s7_c29_n20_c)
    );

    ha ha_s7_c30_n21 (
        .a(stage7_col30[0]),
        .b(stage7_col30[1]),
        .s(ha_s7_c30_n21_s),
        .c_out(ha_s7_c30_n21_c)
    );

    ha ha_s7_c31_n22 (
        .a(stage7_col31[0]),
        .b(stage7_col31[1]),
        .s(ha_s7_c31_n22_s),
        .c_out(ha_s7_c31_n22_c)
    );

    ha ha_s7_c32_n23 (
        .a(stage7_col32[0]),
        .b(stage7_col32[1]),
        .s(ha_s7_c32_n23_s),
        .c_out(ha_s7_c32_n23_c)
    );

    ha ha_s7_c33_n24 (
        .a(stage7_col33[0]),
        .b(stage7_col33[1]),
        .s(ha_s7_c33_n24_s),
        .c_out(ha_s7_c33_n24_c)
    );

    ha ha_s7_c34_n25 (
        .a(stage7_col34[0]),
        .b(stage7_col34[1]),
        .s(ha_s7_c34_n25_s),
        .c_out(ha_s7_c34_n25_c)
    );

    ha ha_s7_c35_n26 (
        .a(stage7_col35[0]),
        .b(stage7_col35[1]),
        .s(ha_s7_c35_n26_s),
        .c_out(ha_s7_c35_n26_c)
    );

    ha ha_s7_c36_n27 (
        .a(stage7_col36[0]),
        .b(stage7_col36[1]),
        .s(ha_s7_c36_n27_s),
        .c_out(ha_s7_c36_n27_c)
    );

    ha ha_s7_c37_n28 (
        .a(stage7_col37[0]),
        .b(stage7_col37[1]),
        .s(ha_s7_c37_n28_s),
        .c_out(ha_s7_c37_n28_c)
    );

    ha ha_s7_c38_n29 (
        .a(stage7_col38[0]),
        .b(stage7_col38[1]),
        .s(ha_s7_c38_n29_s),
        .c_out(ha_s7_c38_n29_c)
    );

    ha ha_s7_c39_n30 (
        .a(stage7_col39[0]),
        .b(stage7_col39[1]),
        .s(ha_s7_c39_n30_s),
        .c_out(ha_s7_c39_n30_c)
    );

    ha ha_s7_c40_n31 (
        .a(stage7_col40[0]),
        .b(stage7_col40[1]),
        .s(ha_s7_c40_n31_s),
        .c_out(ha_s7_c40_n31_c)
    );

    ha ha_s7_c41_n32 (
        .a(stage7_col41[0]),
        .b(stage7_col41[1]),
        .s(ha_s7_c41_n32_s),
        .c_out(ha_s7_c41_n32_c)
    );

    ha ha_s7_c42_n33 (
        .a(stage7_col42[0]),
        .b(stage7_col42[1]),
        .s(ha_s7_c42_n33_s),
        .c_out(ha_s7_c42_n33_c)
    );

    ha ha_s7_c43_n34 (
        .a(stage7_col43[0]),
        .b(stage7_col43[1]),
        .s(ha_s7_c43_n34_s),
        .c_out(ha_s7_c43_n34_c)
    );

    ha ha_s7_c44_n35 (
        .a(stage7_col44[0]),
        .b(stage7_col44[1]),
        .s(ha_s7_c44_n35_s),
        .c_out(ha_s7_c44_n35_c)
    );

    ha ha_s7_c45_n36 (
        .a(stage7_col45[0]),
        .b(stage7_col45[1]),
        .s(ha_s7_c45_n36_s),
        .c_out(ha_s7_c45_n36_c)
    );

    ha ha_s7_c46_n37 (
        .a(stage7_col46[0]),
        .b(stage7_col46[1]),
        .s(ha_s7_c46_n37_s),
        .c_out(ha_s7_c46_n37_c)
    );

    ha ha_s7_c47_n38 (
        .a(stage7_col47[0]),
        .b(stage7_col47[1]),
        .s(ha_s7_c47_n38_s),
        .c_out(ha_s7_c47_n38_c)
    );

    ha ha_s7_c48_n39 (
        .a(stage7_col48[0]),
        .b(stage7_col48[1]),
        .s(ha_s7_c48_n39_s),
        .c_out(ha_s7_c48_n39_c)
    );

    ha ha_s7_c49_n40 (
        .a(stage7_col49[0]),
        .b(stage7_col49[1]),
        .s(ha_s7_c49_n40_s),
        .c_out(ha_s7_c49_n40_c)
    );

    ha ha_s7_c50_n41 (
        .a(stage7_col50[0]),
        .b(stage7_col50[1]),
        .s(ha_s7_c50_n41_s),
        .c_out(ha_s7_c50_n41_c)
    );

    ha ha_s7_c51_n42 (
        .a(stage7_col51[0]),
        .b(stage7_col51[1]),
        .s(ha_s7_c51_n42_s),
        .c_out(ha_s7_c51_n42_c)
    );

    ha ha_s7_c52_n43 (
        .a(stage7_col52[0]),
        .b(stage7_col52[1]),
        .s(ha_s7_c52_n43_s),
        .c_out(ha_s7_c52_n43_c)
    );

    ha ha_s7_c53_n44 (
        .a(stage7_col53[0]),
        .b(stage7_col53[1]),
        .s(ha_s7_c53_n44_s),
        .c_out(ha_s7_c53_n44_c)
    );

    ha ha_s7_c54_n45 (
        .a(stage7_col54[0]),
        .b(stage7_col54[1]),
        .s(ha_s7_c54_n45_s),
        .c_out(ha_s7_c54_n45_c)
    );

    ha ha_s7_c55_n46 (
        .a(stage7_col55[0]),
        .b(stage7_col55[1]),
        .s(ha_s7_c55_n46_s),
        .c_out(ha_s7_c55_n46_c)
    );

    ha ha_s7_c56_n47 (
        .a(stage7_col56[0]),
        .b(stage7_col56[1]),
        .s(ha_s7_c56_n47_s),
        .c_out(ha_s7_c56_n47_c)
    );

    ha ha_s7_c57_n48 (
        .a(stage7_col57[0]),
        .b(stage7_col57[1]),
        .s(ha_s7_c57_n48_s),
        .c_out(ha_s7_c57_n48_c)
    );

    ha ha_s7_c58_n49 (
        .a(stage7_col58[0]),
        .b(stage7_col58[1]),
        .s(ha_s7_c58_n49_s),
        .c_out(ha_s7_c58_n49_c)
    );

    ha ha_s7_c59_n50 (
        .a(stage7_col59[0]),
        .b(stage7_col59[1]),
        .s(ha_s7_c59_n50_s),
        .c_out(ha_s7_c59_n50_c)
    );

    // Map to Stage 8 columns
    generate
        if (PIPE) begin : gen_stage8_pipe
            always_ff @(posedge clk) begin
                if (rst) begin
                    // Reset logic here
                    stage8_col0[0] <= 1'b0;
                    stage8_col1[0] <= 1'b0;
                    stage8_col2[0] <= 1'b0;
                    stage8_col3[0] <= 1'b0;
                    stage8_col4[0] <= 1'b0;
                    stage8_col5[0] <= 1'b0;
                    stage8_col6[0] <= 1'b0;
                    stage8_col7[0] <= 1'b0;
                    stage8_col8[0] <= 1'b0;
                    stage8_col8[1] <= 1'b0;
                    stage8_col9[0] <= 1'b0;
                    stage8_col10[0] <= 1'b0;
                    stage8_col10[1] <= 1'b0;
                    stage8_col11[0] <= 1'b0;
                    stage8_col11[1] <= 1'b0;
                    stage8_col12[0] <= 1'b0;
                    stage8_col12[1] <= 1'b0;
                    stage8_col13[0] <= 1'b0;
                    stage8_col13[1] <= 1'b0;
                    stage8_col14[0] <= 1'b0;
                    stage8_col14[1] <= 1'b0;
                    stage8_col15[0] <= 1'b0;
                    stage8_col15[1] <= 1'b0;
                    stage8_col16[0] <= 1'b0;
                    stage8_col16[1] <= 1'b0;
                    stage8_col17[0] <= 1'b0;
                    stage8_col17[1] <= 1'b0;
                    stage8_col18[0] <= 1'b0;
                    stage8_col18[1] <= 1'b0;
                    stage8_col19[0] <= 1'b0;
                    stage8_col19[1] <= 1'b0;
                    stage8_col20[0] <= 1'b0;
                    stage8_col20[1] <= 1'b0;
                    stage8_col21[0] <= 1'b0;
                    stage8_col21[1] <= 1'b0;
                    stage8_col22[0] <= 1'b0;
                    stage8_col22[1] <= 1'b0;
                    stage8_col23[0] <= 1'b0;
                    stage8_col23[1] <= 1'b0;
                    stage8_col24[0] <= 1'b0;
                    stage8_col24[1] <= 1'b0;
                    stage8_col25[0] <= 1'b0;
                    stage8_col25[1] <= 1'b0;
                    stage8_col26[0] <= 1'b0;
                    stage8_col26[1] <= 1'b0;
                    stage8_col27[0] <= 1'b0;
                    stage8_col27[1] <= 1'b0;
                    stage8_col28[0] <= 1'b0;
                    stage8_col28[1] <= 1'b0;
                    stage8_col29[0] <= 1'b0;
                    stage8_col29[1] <= 1'b0;
                    stage8_col30[0] <= 1'b0;
                    stage8_col30[1] <= 1'b0;
                    stage8_col31[0] <= 1'b0;
                    stage8_col31[1] <= 1'b0;
                    stage8_col32[0] <= 1'b0;
                    stage8_col32[1] <= 1'b0;
                    stage8_col33[0] <= 1'b0;
                    stage8_col33[1] <= 1'b0;
                    stage8_col34[0] <= 1'b0;
                    stage8_col34[1] <= 1'b0;
                    stage8_col35[0] <= 1'b0;
                    stage8_col35[1] <= 1'b0;
                    stage8_col36[0] <= 1'b0;
                    stage8_col36[1] <= 1'b0;
                    stage8_col37[0] <= 1'b0;
                    stage8_col37[1] <= 1'b0;
                    stage8_col38[0] <= 1'b0;
                    stage8_col38[1] <= 1'b0;
                    stage8_col39[0] <= 1'b0;
                    stage8_col39[1] <= 1'b0;
                    stage8_col40[0] <= 1'b0;
                    stage8_col40[1] <= 1'b0;
                    stage8_col41[0] <= 1'b0;
                    stage8_col41[1] <= 1'b0;
                    stage8_col42[0] <= 1'b0;
                    stage8_col42[1] <= 1'b0;
                    stage8_col43[0] <= 1'b0;
                    stage8_col43[1] <= 1'b0;
                    stage8_col44[0] <= 1'b0;
                    stage8_col44[1] <= 1'b0;
                    stage8_col45[0] <= 1'b0;
                    stage8_col45[1] <= 1'b0;
                    stage8_col46[0] <= 1'b0;
                    stage8_col46[1] <= 1'b0;
                    stage8_col47[0] <= 1'b0;
                    stage8_col47[1] <= 1'b0;
                    stage8_col48[0] <= 1'b0;
                    stage8_col48[1] <= 1'b0;
                    stage8_col49[0] <= 1'b0;
                    stage8_col49[1] <= 1'b0;
                    stage8_col50[0] <= 1'b0;
                    stage8_col50[1] <= 1'b0;
                    stage8_col51[0] <= 1'b0;
                    stage8_col51[1] <= 1'b0;
                    stage8_col52[0] <= 1'b0;
                    stage8_col52[1] <= 1'b0;
                    stage8_col53[0] <= 1'b0;
                    stage8_col53[1] <= 1'b0;
                    stage8_col54[0] <= 1'b0;
                    stage8_col54[1] <= 1'b0;
                    stage8_col55[0] <= 1'b0;
                    stage8_col55[1] <= 1'b0;
                    stage8_col56[0] <= 1'b0;
                    stage8_col56[1] <= 1'b0;
                    stage8_col57[0] <= 1'b0;
                    stage8_col57[1] <= 1'b0;
                    stage8_col58[0] <= 1'b0;
                    stage8_col58[1] <= 1'b0;
                    stage8_col59[0] <= 1'b0;
                    stage8_col59[1] <= 1'b0;
                    stage8_col60[0] <= 1'b0;
                    stage8_col60[1] <= 1'b0;
                    stage8_col61[0] <= 1'b0;
                    stage8_col61[1] <= 1'b0;
                    stage8_col62[0] <= 1'b0;
                    stage8_col62[1] <= 1'b0;
                    stage8_col63[0] <= 1'b0;
                    stage8_col63[1] <= 1'b0;
                    stage8_col64[0] <= 1'b0;
                    stage8_col64[1] <= 1'b0;
                    stage8_col65[0] <= 1'b0;
                    stage8_col65[1] <= 1'b0;
                    stage8_col66[0] <= 1'b0;
                    stage8_col66[1] <= 1'b0;
                    stage8_col67[0] <= 1'b0;
                    stage8_col67[1] <= 1'b0;
                    stage8_col68[0] <= 1'b0;
                    stage8_col68[1] <= 1'b0;
                    stage8_col69[0] <= 1'b0;
                    stage8_col69[1] <= 1'b0;
                    stage8_col70[0] <= 1'b0;
                    stage8_col70[1] <= 1'b0;
                    stage8_col71[0] <= 1'b0;
                    stage8_col71[1] <= 1'b0;
                    stage8_col72[0] <= 1'b0;
                    stage8_col72[1] <= 1'b0;
                    stage8_col73[0] <= 1'b0;
                    stage8_col73[1] <= 1'b0;
                    stage8_col74[0] <= 1'b0;
                    stage8_col74[1] <= 1'b0;
                    stage8_col75[0] <= 1'b0;
                    stage8_col75[1] <= 1'b0;
                    stage8_col76[0] <= 1'b0;
                    stage8_col76[1] <= 1'b0;
                    stage8_col77[0] <= 1'b0;
                    stage8_col77[1] <= 1'b0;
                    stage8_col78[0] <= 1'b0;
                    stage8_col78[1] <= 1'b0;
                    stage8_col79[0] <= 1'b0;
                    stage8_col79[1] <= 1'b0;
                    stage8_col80[0] <= 1'b0;
                    stage8_col80[1] <= 1'b0;
                    stage8_col81[0] <= 1'b0;
                    stage8_col81[1] <= 1'b0;
                    stage8_col82[0] <= 1'b0;
                    stage8_col82[1] <= 1'b0;
                    stage8_col83[0] <= 1'b0;
                    stage8_col83[1] <= 1'b0;
                    stage8_col84[0] <= 1'b0;
                    stage8_col84[1] <= 1'b0;
                    stage8_col85[0] <= 1'b0;
                    stage8_col85[1] <= 1'b0;
                    stage8_col86[0] <= 1'b0;
                    stage8_col86[1] <= 1'b0;
                    stage8_col87[0] <= 1'b0;
                    stage8_col87[1] <= 1'b0;
                    stage8_col88[0] <= 1'b0;
                    stage8_col88[1] <= 1'b0;
                    stage8_col89[0] <= 1'b0;
                    stage8_col89[1] <= 1'b0;
                    stage8_col90[0] <= 1'b0;
                    stage8_col90[1] <= 1'b0;
                    stage8_col91[0] <= 1'b0;
                    stage8_col91[1] <= 1'b0;
                    stage8_col92[0] <= 1'b0;
                    stage8_col92[1] <= 1'b0;
                    stage8_col93[0] <= 1'b0;
                    stage8_col93[1] <= 1'b0;
                    stage8_col94[0] <= 1'b0;
                    stage8_col94[1] <= 1'b0;
                    stage8_col95[0] <= 1'b0;
                    stage8_col95[1] <= 1'b0;
                    stage8_col96[0] <= 1'b0;
                    stage8_col96[1] <= 1'b0;
                    stage8_col97[0] <= 1'b0;
                    stage8_col97[1] <= 1'b0;
                    stage8_col98[0] <= 1'b0;
                    stage8_col98[1] <= 1'b0;
                    stage8_col99[0] <= 1'b0;
                    stage8_col99[1] <= 1'b0;
                    stage8_col100[0] <= 1'b0;
                    stage8_col100[1] <= 1'b0;
                    stage8_col101[0] <= 1'b0;
                    stage8_col101[1] <= 1'b0;
                    stage8_col102[0] <= 1'b0;
                    stage8_col102[1] <= 1'b0;
                    stage8_col103[0] <= 1'b0;
                    stage8_col103[1] <= 1'b0;
                    stage8_col104[0] <= 1'b0;
                    stage8_col104[1] <= 1'b0;
                    stage8_col105[0] <= 1'b0;
                    stage8_col105[1] <= 1'b0;
                    stage8_col106[0] <= 1'b0;
                    stage8_col106[1] <= 1'b0;
                    stage8_col107[0] <= 1'b0;
                    stage8_col107[1] <= 1'b0;
                    stage8_col108[0] <= 1'b0;
                    stage8_col108[1] <= 1'b0;
                    stage8_col109[0] <= 1'b0;
                    stage8_col109[1] <= 1'b0;
                    stage8_col110[0] <= 1'b0;
                    stage8_col110[1] <= 1'b0;
                    stage8_col111[0] <= 1'b0;
                    stage8_col111[1] <= 1'b0;
                    stage8_col112[0] <= 1'b0;
                    stage8_col112[1] <= 1'b0;
                    stage8_col113[0] <= 1'b0;
                    stage8_col113[1] <= 1'b0;
                    stage8_col114[0] <= 1'b0;
                    stage8_col114[1] <= 1'b0;
                    stage8_col115[0] <= 1'b0;
                    stage8_col115[1] <= 1'b0;
                    stage8_col116[0] <= 1'b0;
                    stage8_col116[1] <= 1'b0;
                    stage8_col117[0] <= 1'b0;
                    stage8_col117[1] <= 1'b0;
                    stage8_col118[0] <= 1'b0;
                    stage8_col118[1] <= 1'b0;
                    stage8_col119[0] <= 1'b0;
                    stage8_col119[1] <= 1'b0;
                    stage8_col120[0] <= 1'b0;
                    stage8_col120[1] <= 1'b0;
                    stage8_col121[0] <= 1'b0;
                    stage8_col121[1] <= 1'b0;
                    stage8_col122[0] <= 1'b0;
                    stage8_col122[1] <= 1'b0;
                    stage8_col123[0] <= 1'b0;
                    stage8_col123[1] <= 1'b0;
                    stage8_col124[0] <= 1'b0;
                    stage8_col124[1] <= 1'b0;
                    stage8_col125[0] <= 1'b0;
                    stage8_col125[1] <= 1'b0;
                    stage8_col126[0] <= 1'b0;
                    stage8_col126[1] <= 1'b0;
                    stage8_col127[0] <= 1'b0;
                    stage8_col127[1] <= 1'b0;
                    stage8_col127[2] <= 1'b0;
                    stage8_col127[3] <= 1'b0;
                    stage8_col127[4] <= 1'b0;
                    stage8_col127[5] <= 1'b0;
                    stage8_col127[6] <= 1'b0;
                    stage8_col127[7] <= 1'b0;
                    stage8_col127[8] <= 1'b0;
                    stage8_col127[9] <= 1'b0;
                    stage8_col127[10] <= 1'b0;
                    stage8_col127[11] <= 1'b0;
                    stage8_col127[12] <= 1'b0;
                    stage8_col127[13] <= 1'b0;
                    stage8_col127[14] <= 1'b0;
                    stage8_col127[15] <= 1'b0;
                    stage8_col127[16] <= 1'b0;
                    stage8_col127[17] <= 1'b0;
                    stage8_col127[18] <= 1'b0;
                    stage8_col127[19] <= 1'b0;
                    stage8_col127[20] <= 1'b0;
                    stage8_col127[21] <= 1'b0;
                    stage8_col127[22] <= 1'b0;
                    stage8_col127[23] <= 1'b0;
                    stage8_col127[24] <= 1'b0;
                    stage8_col127[25] <= 1'b0;
                    stage8_col127[26] <= 1'b0;
                    stage8_col127[27] <= 1'b0;
                    stage8_col127[28] <= 1'b0;
                    stage8_col127[29] <= 1'b0;
                    stage8_col127[30] <= 1'b0;
                    stage8_col127[31] <= 1'b0;
                    stage8_col127[32] <= 1'b0;
                    stage8_col127[33] <= 1'b0;
                    stage8_col127[34] <= 1'b0;
                    stage8_col127[35] <= 1'b0;
                    stage8_col127[36] <= 1'b0;
                    stage8_col127[37] <= 1'b0;
                    stage8_col127[38] <= 1'b0;
                    stage8_col127[39] <= 1'b0;
                    stage8_col127[40] <= 1'b0;
                    stage8_col127[41] <= 1'b0;
                    stage8_col127[42] <= 1'b0;
                    stage8_col127[43] <= 1'b0;
                    stage8_col127[44] <= 1'b0;
                    stage8_col127[45] <= 1'b0;
                    stage8_col127[46] <= 1'b0;
                    stage8_col127[47] <= 1'b0;
                    stage8_col127[48] <= 1'b0;
                    stage8_col127[49] <= 1'b0;
                    stage8_col127[50] <= 1'b0;
                    stage8_col127[51] <= 1'b0;
                    stage8_col127[52] <= 1'b0;
                    stage8_col127[53] <= 1'b0;
                    stage8_col127[54] <= 1'b0;
                    stage8_col127[55] <= 1'b0;
                    stage8_col127[56] <= 1'b0;
                    stage8_col127[57] <= 1'b0;
                    stage8_col127[58] <= 1'b0;
                    stage8_col127[59] <= 1'b0;
                    stage8_col127[60] <= 1'b0;
                    stage8_col127[61] <= 1'b0;
                    stage8_col127[62] <= 1'b0;
                end else begin
                    // Normal operation logic here
                    stage8_col0[0] <= stage7_col0[0];
                    stage8_col1[0] <= stage7_col1[0];
                    stage8_col2[0] <= stage7_col2[0];
                    stage8_col3[0] <= stage7_col3[0];
                    stage8_col4[0] <= stage7_col4[0];
                    stage8_col5[0] <= stage7_col5[0];
                    stage8_col6[0] <= stage7_col6[0];
                    stage8_col7[0] <= ha_s7_c7_n0_s;
                    stage8_col8[0] <= ha_s7_c7_n0_c;
                    stage8_col8[1] <= stage7_col8[0];
                    stage8_col9[0] <= fa_s7_c9_n0_s;
                    stage8_col10[0] <= fa_s7_c9_n0_c;
                    stage8_col10[1] <= ha_s7_c10_n1_s;
                    stage8_col11[0] <= ha_s7_c10_n1_c;
                    stage8_col11[1] <= ha_s7_c11_n2_s;
                    stage8_col12[0] <= ha_s7_c11_n2_c;
                    stage8_col12[1] <= ha_s7_c12_n3_s;
                    stage8_col13[0] <= ha_s7_c12_n3_c;
                    stage8_col13[1] <= ha_s7_c13_n4_s;
                    stage8_col14[0] <= ha_s7_c13_n4_c;
                    stage8_col14[1] <= ha_s7_c14_n5_s;
                    stage8_col15[0] <= ha_s7_c14_n5_c;
                    stage8_col15[1] <= ha_s7_c15_n6_s;
                    stage8_col16[0] <= ha_s7_c15_n6_c;
                    stage8_col16[1] <= ha_s7_c16_n7_s;
                    stage8_col17[0] <= ha_s7_c16_n7_c;
                    stage8_col17[1] <= ha_s7_c17_n8_s;
                    stage8_col18[0] <= ha_s7_c17_n8_c;
                    stage8_col18[1] <= ha_s7_c18_n9_s;
                    stage8_col19[0] <= ha_s7_c18_n9_c;
                    stage8_col19[1] <= ha_s7_c19_n10_s;
                    stage8_col20[0] <= ha_s7_c19_n10_c;
                    stage8_col20[1] <= ha_s7_c20_n11_s;
                    stage8_col21[0] <= ha_s7_c20_n11_c;
                    stage8_col21[1] <= ha_s7_c21_n12_s;
                    stage8_col22[0] <= ha_s7_c21_n12_c;
                    stage8_col22[1] <= ha_s7_c22_n13_s;
                    stage8_col23[0] <= ha_s7_c22_n13_c;
                    stage8_col23[1] <= ha_s7_c23_n14_s;
                    stage8_col24[0] <= ha_s7_c23_n14_c;
                    stage8_col24[1] <= ha_s7_c24_n15_s;
                    stage8_col25[0] <= ha_s7_c24_n15_c;
                    stage8_col25[1] <= ha_s7_c25_n16_s;
                    stage8_col26[0] <= ha_s7_c25_n16_c;
                    stage8_col26[1] <= ha_s7_c26_n17_s;
                    stage8_col27[0] <= ha_s7_c26_n17_c;
                    stage8_col27[1] <= ha_s7_c27_n18_s;
                    stage8_col28[0] <= ha_s7_c27_n18_c;
                    stage8_col28[1] <= ha_s7_c28_n19_s;
                    stage8_col29[0] <= ha_s7_c28_n19_c;
                    stage8_col29[1] <= ha_s7_c29_n20_s;
                    stage8_col30[0] <= ha_s7_c29_n20_c;
                    stage8_col30[1] <= ha_s7_c30_n21_s;
                    stage8_col31[0] <= ha_s7_c30_n21_c;
                    stage8_col31[1] <= ha_s7_c31_n22_s;
                    stage8_col32[0] <= ha_s7_c31_n22_c;
                    stage8_col32[1] <= ha_s7_c32_n23_s;
                    stage8_col33[0] <= ha_s7_c32_n23_c;
                    stage8_col33[1] <= ha_s7_c33_n24_s;
                    stage8_col34[0] <= ha_s7_c33_n24_c;
                    stage8_col34[1] <= ha_s7_c34_n25_s;
                    stage8_col35[0] <= ha_s7_c34_n25_c;
                    stage8_col35[1] <= ha_s7_c35_n26_s;
                    stage8_col36[0] <= ha_s7_c35_n26_c;
                    stage8_col36[1] <= ha_s7_c36_n27_s;
                    stage8_col37[0] <= ha_s7_c36_n27_c;
                    stage8_col37[1] <= ha_s7_c37_n28_s;
                    stage8_col38[0] <= ha_s7_c37_n28_c;
                    stage8_col38[1] <= ha_s7_c38_n29_s;
                    stage8_col39[0] <= ha_s7_c38_n29_c;
                    stage8_col39[1] <= ha_s7_c39_n30_s;
                    stage8_col40[0] <= ha_s7_c39_n30_c;
                    stage8_col40[1] <= ha_s7_c40_n31_s;
                    stage8_col41[0] <= ha_s7_c40_n31_c;
                    stage8_col41[1] <= ha_s7_c41_n32_s;
                    stage8_col42[0] <= ha_s7_c41_n32_c;
                    stage8_col42[1] <= ha_s7_c42_n33_s;
                    stage8_col43[0] <= ha_s7_c42_n33_c;
                    stage8_col43[1] <= ha_s7_c43_n34_s;
                    stage8_col44[0] <= ha_s7_c43_n34_c;
                    stage8_col44[1] <= ha_s7_c44_n35_s;
                    stage8_col45[0] <= ha_s7_c44_n35_c;
                    stage8_col45[1] <= ha_s7_c45_n36_s;
                    stage8_col46[0] <= ha_s7_c45_n36_c;
                    stage8_col46[1] <= ha_s7_c46_n37_s;
                    stage8_col47[0] <= ha_s7_c46_n37_c;
                    stage8_col47[1] <= ha_s7_c47_n38_s;
                    stage8_col48[0] <= ha_s7_c47_n38_c;
                    stage8_col48[1] <= ha_s7_c48_n39_s;
                    stage8_col49[0] <= ha_s7_c48_n39_c;
                    stage8_col49[1] <= ha_s7_c49_n40_s;
                    stage8_col50[0] <= ha_s7_c49_n40_c;
                    stage8_col50[1] <= ha_s7_c50_n41_s;
                    stage8_col51[0] <= ha_s7_c50_n41_c;
                    stage8_col51[1] <= ha_s7_c51_n42_s;
                    stage8_col52[0] <= ha_s7_c51_n42_c;
                    stage8_col52[1] <= ha_s7_c52_n43_s;
                    stage8_col53[0] <= ha_s7_c52_n43_c;
                    stage8_col53[1] <= ha_s7_c53_n44_s;
                    stage8_col54[0] <= ha_s7_c53_n44_c;
                    stage8_col54[1] <= ha_s7_c54_n45_s;
                    stage8_col55[0] <= ha_s7_c54_n45_c;
                    stage8_col55[1] <= ha_s7_c55_n46_s;
                    stage8_col56[0] <= ha_s7_c55_n46_c;
                    stage8_col56[1] <= ha_s7_c56_n47_s;
                    stage8_col57[0] <= ha_s7_c56_n47_c;
                    stage8_col57[1] <= ha_s7_c57_n48_s;
                    stage8_col58[0] <= ha_s7_c57_n48_c;
                    stage8_col58[1] <= ha_s7_c58_n49_s;
                    stage8_col59[0] <= ha_s7_c58_n49_c;
                    stage8_col59[1] <= ha_s7_c59_n50_s;
                    stage8_col60[0] <= ha_s7_c59_n50_c;
                    stage8_col60[1] <= fa_s7_c60_n1_s;
                    stage8_col61[0] <= fa_s7_c60_n1_c;
                    stage8_col61[1] <= fa_s7_c61_n2_s;
                    stage8_col62[0] <= fa_s7_c61_n2_c;
                    stage8_col62[1] <= fa_s7_c62_n3_s;
                    stage8_col63[0] <= fa_s7_c62_n3_c;
                    stage8_col63[1] <= fa_s7_c63_n4_s;
                    stage8_col64[0] <= fa_s7_c63_n4_c;
                    stage8_col64[1] <= fa_s7_c64_n5_s;
                    stage8_col65[0] <= fa_s7_c64_n5_c;
                    stage8_col65[1] <= fa_s7_c65_n6_s;
                    stage8_col66[0] <= fa_s7_c65_n6_c;
                    stage8_col66[1] <= fa_s7_c66_n7_s;
                    stage8_col67[0] <= fa_s7_c66_n7_c;
                    stage8_col67[1] <= fa_s7_c67_n8_s;
                    stage8_col68[0] <= fa_s7_c67_n8_c;
                    stage8_col68[1] <= fa_s7_c68_n9_s;
                    stage8_col69[0] <= fa_s7_c68_n9_c;
                    stage8_col69[1] <= fa_s7_c69_n10_s;
                    stage8_col70[0] <= fa_s7_c69_n10_c;
                    stage8_col70[1] <= fa_s7_c70_n11_s;
                    stage8_col71[0] <= fa_s7_c70_n11_c;
                    stage8_col71[1] <= fa_s7_c71_n12_s;
                    stage8_col72[0] <= fa_s7_c71_n12_c;
                    stage8_col72[1] <= fa_s7_c72_n13_s;
                    stage8_col73[0] <= fa_s7_c72_n13_c;
                    stage8_col73[1] <= fa_s7_c73_n14_s;
                    stage8_col74[0] <= fa_s7_c73_n14_c;
                    stage8_col74[1] <= fa_s7_c74_n15_s;
                    stage8_col75[0] <= fa_s7_c74_n15_c;
                    stage8_col75[1] <= fa_s7_c75_n16_s;
                    stage8_col76[0] <= fa_s7_c75_n16_c;
                    stage8_col76[1] <= fa_s7_c76_n17_s;
                    stage8_col77[0] <= fa_s7_c76_n17_c;
                    stage8_col77[1] <= fa_s7_c77_n18_s;
                    stage8_col78[0] <= fa_s7_c77_n18_c;
                    stage8_col78[1] <= fa_s7_c78_n19_s;
                    stage8_col79[0] <= fa_s7_c78_n19_c;
                    stage8_col79[1] <= fa_s7_c79_n20_s;
                    stage8_col80[0] <= fa_s7_c79_n20_c;
                    stage8_col80[1] <= fa_s7_c80_n21_s;
                    stage8_col81[0] <= fa_s7_c80_n21_c;
                    stage8_col81[1] <= fa_s7_c81_n22_s;
                    stage8_col82[0] <= fa_s7_c81_n22_c;
                    stage8_col82[1] <= fa_s7_c82_n23_s;
                    stage8_col83[0] <= fa_s7_c82_n23_c;
                    stage8_col83[1] <= fa_s7_c83_n24_s;
                    stage8_col84[0] <= fa_s7_c83_n24_c;
                    stage8_col84[1] <= fa_s7_c84_n25_s;
                    stage8_col85[0] <= fa_s7_c84_n25_c;
                    stage8_col85[1] <= fa_s7_c85_n26_s;
                    stage8_col86[0] <= fa_s7_c85_n26_c;
                    stage8_col86[1] <= fa_s7_c86_n27_s;
                    stage8_col87[0] <= fa_s7_c86_n27_c;
                    stage8_col87[1] <= fa_s7_c87_n28_s;
                    stage8_col88[0] <= fa_s7_c87_n28_c;
                    stage8_col88[1] <= fa_s7_c88_n29_s;
                    stage8_col89[0] <= fa_s7_c88_n29_c;
                    stage8_col89[1] <= fa_s7_c89_n30_s;
                    stage8_col90[0] <= fa_s7_c89_n30_c;
                    stage8_col90[1] <= fa_s7_c90_n31_s;
                    stage8_col91[0] <= fa_s7_c90_n31_c;
                    stage8_col91[1] <= fa_s7_c91_n32_s;
                    stage8_col92[0] <= fa_s7_c91_n32_c;
                    stage8_col92[1] <= fa_s7_c92_n33_s;
                    stage8_col93[0] <= fa_s7_c92_n33_c;
                    stage8_col93[1] <= fa_s7_c93_n34_s;
                    stage8_col94[0] <= fa_s7_c93_n34_c;
                    stage8_col94[1] <= fa_s7_c94_n35_s;
                    stage8_col95[0] <= fa_s7_c94_n35_c;
                    stage8_col95[1] <= fa_s7_c95_n36_s;
                    stage8_col96[0] <= fa_s7_c95_n36_c;
                    stage8_col96[1] <= fa_s7_c96_n37_s;
                    stage8_col97[0] <= fa_s7_c96_n37_c;
                    stage8_col97[1] <= fa_s7_c97_n38_s;
                    stage8_col98[0] <= fa_s7_c97_n38_c;
                    stage8_col98[1] <= fa_s7_c98_n39_s;
                    stage8_col99[0] <= fa_s7_c98_n39_c;
                    stage8_col99[1] <= fa_s7_c99_n40_s;
                    stage8_col100[0] <= fa_s7_c99_n40_c;
                    stage8_col100[1] <= fa_s7_c100_n41_s;
                    stage8_col101[0] <= fa_s7_c100_n41_c;
                    stage8_col101[1] <= fa_s7_c101_n42_s;
                    stage8_col102[0] <= fa_s7_c101_n42_c;
                    stage8_col102[1] <= fa_s7_c102_n43_s;
                    stage8_col103[0] <= fa_s7_c102_n43_c;
                    stage8_col103[1] <= fa_s7_c103_n44_s;
                    stage8_col104[0] <= fa_s7_c103_n44_c;
                    stage8_col104[1] <= fa_s7_c104_n45_s;
                    stage8_col105[0] <= fa_s7_c104_n45_c;
                    stage8_col105[1] <= fa_s7_c105_n46_s;
                    stage8_col106[0] <= fa_s7_c105_n46_c;
                    stage8_col106[1] <= fa_s7_c106_n47_s;
                    stage8_col107[0] <= fa_s7_c106_n47_c;
                    stage8_col107[1] <= fa_s7_c107_n48_s;
                    stage8_col108[0] <= fa_s7_c107_n48_c;
                    stage8_col108[1] <= fa_s7_c108_n49_s;
                    stage8_col109[0] <= fa_s7_c108_n49_c;
                    stage8_col109[1] <= fa_s7_c109_n50_s;
                    stage8_col110[0] <= fa_s7_c109_n50_c;
                    stage8_col110[1] <= fa_s7_c110_n51_s;
                    stage8_col111[0] <= fa_s7_c110_n51_c;
                    stage8_col111[1] <= fa_s7_c111_n52_s;
                    stage8_col112[0] <= fa_s7_c111_n52_c;
                    stage8_col112[1] <= fa_s7_c112_n53_s;
                    stage8_col113[0] <= fa_s7_c112_n53_c;
                    stage8_col113[1] <= fa_s7_c113_n54_s;
                    stage8_col114[0] <= fa_s7_c113_n54_c;
                    stage8_col114[1] <= fa_s7_c114_n55_s;
                    stage8_col115[0] <= fa_s7_c114_n55_c;
                    stage8_col115[1] <= fa_s7_c115_n56_s;
                    stage8_col116[0] <= fa_s7_c115_n56_c;
                    stage8_col116[1] <= fa_s7_c116_n57_s;
                    stage8_col117[0] <= fa_s7_c116_n57_c;
                    stage8_col117[1] <= fa_s7_c117_n58_s;
                    stage8_col118[0] <= fa_s7_c117_n58_c;
                    stage8_col118[1] <= fa_s7_c118_n59_s;
                    stage8_col119[0] <= fa_s7_c118_n59_c;
                    stage8_col119[1] <= fa_s7_c119_n60_s;
                    stage8_col120[0] <= fa_s7_c119_n60_c;
                    stage8_col120[1] <= fa_s7_c120_n61_s;
                    stage8_col121[0] <= fa_s7_c120_n61_c;
                    stage8_col121[1] <= fa_s7_c121_n62_s;
                    stage8_col122[0] <= fa_s7_c121_n62_c;
                    stage8_col122[1] <= fa_s7_c122_n63_s;
                    stage8_col123[0] <= fa_s7_c122_n63_c;
                    stage8_col123[1] <= fa_s7_c123_n64_s;
                    stage8_col124[0] <= fa_s7_c123_n64_c;
                    stage8_col124[1] <= fa_s7_c124_n65_s;
                    stage8_col125[0] <= fa_s7_c124_n65_c;
                    stage8_col125[1] <= fa_s7_c125_n66_s;
                    stage8_col126[0] <= fa_s7_c125_n66_c;
                    stage8_col126[1] <= fa_s7_c126_n67_s;
                    stage8_col127[0] <= fa_s7_c126_n67_c;
                    stage8_col127[1] <= stage7_col127[0];
                    stage8_col127[2] <= stage7_col127[1];
                    stage8_col127[3] <= stage7_col127[2];
                    stage8_col127[4] <= stage7_col127[3];
                    stage8_col127[5] <= stage7_col127[4];
                    stage8_col127[6] <= stage7_col127[5];
                    stage8_col127[7] <= stage7_col127[6];
                    stage8_col127[8] <= stage7_col127[7];
                    stage8_col127[9] <= stage7_col127[8];
                    stage8_col127[10] <= stage7_col127[9];
                    stage8_col127[11] <= stage7_col127[10];
                    stage8_col127[12] <= stage7_col127[11];
                    stage8_col127[13] <= stage7_col127[12];
                    stage8_col127[14] <= stage7_col127[13];
                    stage8_col127[15] <= stage7_col127[14];
                    stage8_col127[16] <= stage7_col127[15];
                    stage8_col127[17] <= stage7_col127[16];
                    stage8_col127[18] <= stage7_col127[17];
                    stage8_col127[19] <= stage7_col127[18];
                    stage8_col127[20] <= stage7_col127[19];
                    stage8_col127[21] <= stage7_col127[20];
                    stage8_col127[22] <= stage7_col127[21];
                    stage8_col127[23] <= stage7_col127[22];
                    stage8_col127[24] <= stage7_col127[23];
                    stage8_col127[25] <= stage7_col127[24];
                    stage8_col127[26] <= stage7_col127[25];
                    stage8_col127[27] <= stage7_col127[26];
                    stage8_col127[28] <= stage7_col127[27];
                    stage8_col127[29] <= stage7_col127[28];
                    stage8_col127[30] <= stage7_col127[29];
                    stage8_col127[31] <= stage7_col127[30];
                    stage8_col127[32] <= stage7_col127[30];
                    stage8_col127[33] <= stage7_col127[30];
                    stage8_col127[34] <= stage7_col127[30];
                    stage8_col127[35] <= stage7_col127[30];
                    stage8_col127[36] <= stage7_col127[30];
                    stage8_col127[37] <= stage7_col127[30];
                    stage8_col127[38] <= stage7_col127[30];
                    stage8_col127[39] <= stage7_col127[30];
                    stage8_col127[40] <= stage7_col127[30];
                    stage8_col127[41] <= stage7_col127[30];
                    stage8_col127[42] <= stage7_col127[30];
                    stage8_col127[43] <= stage7_col127[30];
                    stage8_col127[44] <= stage7_col127[30];
                    stage8_col127[45] <= stage7_col127[30];
                    stage8_col127[46] <= stage7_col127[30];
                    stage8_col127[47] <= stage7_col127[30];
                    stage8_col127[48] <= stage7_col127[30];
                    stage8_col127[49] <= stage7_col127[30];
                    stage8_col127[50] <= stage7_col127[30];
                    stage8_col127[51] <= stage7_col127[30];
                    stage8_col127[52] <= stage7_col127[30];
                    stage8_col127[53] <= stage7_col127[30];
                    stage8_col127[54] <= stage7_col127[30];
                    stage8_col127[55] <= stage7_col127[30];
                    stage8_col127[56] <= stage7_col127[30];
                    stage8_col127[57] <= stage7_col127[30];
                    stage8_col127[58] <= stage7_col127[30];
                    stage8_col127[59] <= stage7_col127[30];
                    stage8_col127[60] <= stage7_col127[30];
                    stage8_col127[61] <= stage7_col127[30];
                    stage8_col127[62] <= stage7_col127[30];
                end
            end
        end else begin : gen_stage8_no_pipe
            // Combinational assignment
            always_comb begin
                stage8_col0[0] = stage7_col0[0];
                stage8_col1[0] = stage7_col1[0];
                stage8_col2[0] = stage7_col2[0];
                stage8_col3[0] = stage7_col3[0];
                stage8_col4[0] = stage7_col4[0];
                stage8_col5[0] = stage7_col5[0];
                stage8_col6[0] = stage7_col6[0];
                stage8_col7[0] = ha_s7_c7_n0_s;
                stage8_col8[0] = ha_s7_c7_n0_c;
                stage8_col8[1] = stage7_col8[0];
                stage8_col9[0] = fa_s7_c9_n0_s;
                stage8_col10[0] = fa_s7_c9_n0_c;
                stage8_col10[1] = ha_s7_c10_n1_s;
                stage8_col11[0] = ha_s7_c10_n1_c;
                stage8_col11[1] = ha_s7_c11_n2_s;
                stage8_col12[0] = ha_s7_c11_n2_c;
                stage8_col12[1] = ha_s7_c12_n3_s;
                stage8_col13[0] = ha_s7_c12_n3_c;
                stage8_col13[1] = ha_s7_c13_n4_s;
                stage8_col14[0] = ha_s7_c13_n4_c;
                stage8_col14[1] = ha_s7_c14_n5_s;
                stage8_col15[0] = ha_s7_c14_n5_c;
                stage8_col15[1] = ha_s7_c15_n6_s;
                stage8_col16[0] = ha_s7_c15_n6_c;
                stage8_col16[1] = ha_s7_c16_n7_s;
                stage8_col17[0] = ha_s7_c16_n7_c;
                stage8_col17[1] = ha_s7_c17_n8_s;
                stage8_col18[0] = ha_s7_c17_n8_c;
                stage8_col18[1] = ha_s7_c18_n9_s;
                stage8_col19[0] = ha_s7_c18_n9_c;
                stage8_col19[1] = ha_s7_c19_n10_s;
                stage8_col20[0] = ha_s7_c19_n10_c;
                stage8_col20[1] = ha_s7_c20_n11_s;
                stage8_col21[0] = ha_s7_c20_n11_c;
                stage8_col21[1] = ha_s7_c21_n12_s;
                stage8_col22[0] = ha_s7_c21_n12_c;
                stage8_col22[1] = ha_s7_c22_n13_s;
                stage8_col23[0] = ha_s7_c22_n13_c;
                stage8_col23[1] = ha_s7_c23_n14_s;
                stage8_col24[0] = ha_s7_c23_n14_c;
                stage8_col24[1] = ha_s7_c24_n15_s;
                stage8_col25[0] = ha_s7_c24_n15_c;
                stage8_col25[1] = ha_s7_c25_n16_s;
                stage8_col26[0] = ha_s7_c25_n16_c;
                stage8_col26[1] = ha_s7_c26_n17_s;
                stage8_col27[0] = ha_s7_c26_n17_c;
                stage8_col27[1] = ha_s7_c27_n18_s;
                stage8_col28[0] = ha_s7_c27_n18_c;
                stage8_col28[1] = ha_s7_c28_n19_s;
                stage8_col29[0] = ha_s7_c28_n19_c;
                stage8_col29[1] = ha_s7_c29_n20_s;
                stage8_col30[0] = ha_s7_c29_n20_c;
                stage8_col30[1] = ha_s7_c30_n21_s;
                stage8_col31[0] = ha_s7_c30_n21_c;
                stage8_col31[1] = ha_s7_c31_n22_s;
                stage8_col32[0] = ha_s7_c31_n22_c;
                stage8_col32[1] = ha_s7_c32_n23_s;
                stage8_col33[0] = ha_s7_c32_n23_c;
                stage8_col33[1] = ha_s7_c33_n24_s;
                stage8_col34[0] = ha_s7_c33_n24_c;
                stage8_col34[1] = ha_s7_c34_n25_s;
                stage8_col35[0] = ha_s7_c34_n25_c;
                stage8_col35[1] = ha_s7_c35_n26_s;
                stage8_col36[0] = ha_s7_c35_n26_c;
                stage8_col36[1] = ha_s7_c36_n27_s;
                stage8_col37[0] = ha_s7_c36_n27_c;
                stage8_col37[1] = ha_s7_c37_n28_s;
                stage8_col38[0] = ha_s7_c37_n28_c;
                stage8_col38[1] = ha_s7_c38_n29_s;
                stage8_col39[0] = ha_s7_c38_n29_c;
                stage8_col39[1] = ha_s7_c39_n30_s;
                stage8_col40[0] = ha_s7_c39_n30_c;
                stage8_col40[1] = ha_s7_c40_n31_s;
                stage8_col41[0] = ha_s7_c40_n31_c;
                stage8_col41[1] = ha_s7_c41_n32_s;
                stage8_col42[0] = ha_s7_c41_n32_c;
                stage8_col42[1] = ha_s7_c42_n33_s;
                stage8_col43[0] = ha_s7_c42_n33_c;
                stage8_col43[1] = ha_s7_c43_n34_s;
                stage8_col44[0] = ha_s7_c43_n34_c;
                stage8_col44[1] = ha_s7_c44_n35_s;
                stage8_col45[0] = ha_s7_c44_n35_c;
                stage8_col45[1] = ha_s7_c45_n36_s;
                stage8_col46[0] = ha_s7_c45_n36_c;
                stage8_col46[1] = ha_s7_c46_n37_s;
                stage8_col47[0] = ha_s7_c46_n37_c;
                stage8_col47[1] = ha_s7_c47_n38_s;
                stage8_col48[0] = ha_s7_c47_n38_c;
                stage8_col48[1] = ha_s7_c48_n39_s;
                stage8_col49[0] = ha_s7_c48_n39_c;
                stage8_col49[1] = ha_s7_c49_n40_s;
                stage8_col50[0] = ha_s7_c49_n40_c;
                stage8_col50[1] = ha_s7_c50_n41_s;
                stage8_col51[0] = ha_s7_c50_n41_c;
                stage8_col51[1] = ha_s7_c51_n42_s;
                stage8_col52[0] = ha_s7_c51_n42_c;
                stage8_col52[1] = ha_s7_c52_n43_s;
                stage8_col53[0] = ha_s7_c52_n43_c;
                stage8_col53[1] = ha_s7_c53_n44_s;
                stage8_col54[0] = ha_s7_c53_n44_c;
                stage8_col54[1] = ha_s7_c54_n45_s;
                stage8_col55[0] = ha_s7_c54_n45_c;
                stage8_col55[1] = ha_s7_c55_n46_s;
                stage8_col56[0] = ha_s7_c55_n46_c;
                stage8_col56[1] = ha_s7_c56_n47_s;
                stage8_col57[0] = ha_s7_c56_n47_c;
                stage8_col57[1] = ha_s7_c57_n48_s;
                stage8_col58[0] = ha_s7_c57_n48_c;
                stage8_col58[1] = ha_s7_c58_n49_s;
                stage8_col59[0] = ha_s7_c58_n49_c;
                stage8_col59[1] = ha_s7_c59_n50_s;
                stage8_col60[0] = ha_s7_c59_n50_c;
                stage8_col60[1] = fa_s7_c60_n1_s;
                stage8_col61[0] = fa_s7_c60_n1_c;
                stage8_col61[1] = fa_s7_c61_n2_s;
                stage8_col62[0] = fa_s7_c61_n2_c;
                stage8_col62[1] = fa_s7_c62_n3_s;
                stage8_col63[0] = fa_s7_c62_n3_c;
                stage8_col63[1] = fa_s7_c63_n4_s;
                stage8_col64[0] = fa_s7_c63_n4_c;
                stage8_col64[1] = fa_s7_c64_n5_s;
                stage8_col65[0] = fa_s7_c64_n5_c;
                stage8_col65[1] = fa_s7_c65_n6_s;
                stage8_col66[0] = fa_s7_c65_n6_c;
                stage8_col66[1] = fa_s7_c66_n7_s;
                stage8_col67[0] = fa_s7_c66_n7_c;
                stage8_col67[1] = fa_s7_c67_n8_s;
                stage8_col68[0] = fa_s7_c67_n8_c;
                stage8_col68[1] = fa_s7_c68_n9_s;
                stage8_col69[0] = fa_s7_c68_n9_c;
                stage8_col69[1] = fa_s7_c69_n10_s;
                stage8_col70[0] = fa_s7_c69_n10_c;
                stage8_col70[1] = fa_s7_c70_n11_s;
                stage8_col71[0] = fa_s7_c70_n11_c;
                stage8_col71[1] = fa_s7_c71_n12_s;
                stage8_col72[0] = fa_s7_c71_n12_c;
                stage8_col72[1] = fa_s7_c72_n13_s;
                stage8_col73[0] = fa_s7_c72_n13_c;
                stage8_col73[1] = fa_s7_c73_n14_s;
                stage8_col74[0] = fa_s7_c73_n14_c;
                stage8_col74[1] = fa_s7_c74_n15_s;
                stage8_col75[0] = fa_s7_c74_n15_c;
                stage8_col75[1] = fa_s7_c75_n16_s;
                stage8_col76[0] = fa_s7_c75_n16_c;
                stage8_col76[1] = fa_s7_c76_n17_s;
                stage8_col77[0] = fa_s7_c76_n17_c;
                stage8_col77[1] = fa_s7_c77_n18_s;
                stage8_col78[0] = fa_s7_c77_n18_c;
                stage8_col78[1] = fa_s7_c78_n19_s;
                stage8_col79[0] = fa_s7_c78_n19_c;
                stage8_col79[1] = fa_s7_c79_n20_s;
                stage8_col80[0] = fa_s7_c79_n20_c;
                stage8_col80[1] = fa_s7_c80_n21_s;
                stage8_col81[0] = fa_s7_c80_n21_c;
                stage8_col81[1] = fa_s7_c81_n22_s;
                stage8_col82[0] = fa_s7_c81_n22_c;
                stage8_col82[1] = fa_s7_c82_n23_s;
                stage8_col83[0] = fa_s7_c82_n23_c;
                stage8_col83[1] = fa_s7_c83_n24_s;
                stage8_col84[0] = fa_s7_c83_n24_c;
                stage8_col84[1] = fa_s7_c84_n25_s;
                stage8_col85[0] = fa_s7_c84_n25_c;
                stage8_col85[1] = fa_s7_c85_n26_s;
                stage8_col86[0] = fa_s7_c85_n26_c;
                stage8_col86[1] = fa_s7_c86_n27_s;
                stage8_col87[0] = fa_s7_c86_n27_c;
                stage8_col87[1] = fa_s7_c87_n28_s;
                stage8_col88[0] = fa_s7_c87_n28_c;
                stage8_col88[1] = fa_s7_c88_n29_s;
                stage8_col89[0] = fa_s7_c88_n29_c;
                stage8_col89[1] = fa_s7_c89_n30_s;
                stage8_col90[0] = fa_s7_c89_n30_c;
                stage8_col90[1] = fa_s7_c90_n31_s;
                stage8_col91[0] = fa_s7_c90_n31_c;
                stage8_col91[1] = fa_s7_c91_n32_s;
                stage8_col92[0] = fa_s7_c91_n32_c;
                stage8_col92[1] = fa_s7_c92_n33_s;
                stage8_col93[0] = fa_s7_c92_n33_c;
                stage8_col93[1] = fa_s7_c93_n34_s;
                stage8_col94[0] = fa_s7_c93_n34_c;
                stage8_col94[1] = fa_s7_c94_n35_s;
                stage8_col95[0] = fa_s7_c94_n35_c;
                stage8_col95[1] = fa_s7_c95_n36_s;
                stage8_col96[0] = fa_s7_c95_n36_c;
                stage8_col96[1] = fa_s7_c96_n37_s;
                stage8_col97[0] = fa_s7_c96_n37_c;
                stage8_col97[1] = fa_s7_c97_n38_s;
                stage8_col98[0] = fa_s7_c97_n38_c;
                stage8_col98[1] = fa_s7_c98_n39_s;
                stage8_col99[0] = fa_s7_c98_n39_c;
                stage8_col99[1] = fa_s7_c99_n40_s;
                stage8_col100[0] = fa_s7_c99_n40_c;
                stage8_col100[1] = fa_s7_c100_n41_s;
                stage8_col101[0] = fa_s7_c100_n41_c;
                stage8_col101[1] = fa_s7_c101_n42_s;
                stage8_col102[0] = fa_s7_c101_n42_c;
                stage8_col102[1] = fa_s7_c102_n43_s;
                stage8_col103[0] = fa_s7_c102_n43_c;
                stage8_col103[1] = fa_s7_c103_n44_s;
                stage8_col104[0] = fa_s7_c103_n44_c;
                stage8_col104[1] = fa_s7_c104_n45_s;
                stage8_col105[0] = fa_s7_c104_n45_c;
                stage8_col105[1] = fa_s7_c105_n46_s;
                stage8_col106[0] = fa_s7_c105_n46_c;
                stage8_col106[1] = fa_s7_c106_n47_s;
                stage8_col107[0] = fa_s7_c106_n47_c;
                stage8_col107[1] = fa_s7_c107_n48_s;
                stage8_col108[0] = fa_s7_c107_n48_c;
                stage8_col108[1] = fa_s7_c108_n49_s;
                stage8_col109[0] = fa_s7_c108_n49_c;
                stage8_col109[1] = fa_s7_c109_n50_s;
                stage8_col110[0] = fa_s7_c109_n50_c;
                stage8_col110[1] = fa_s7_c110_n51_s;
                stage8_col111[0] = fa_s7_c110_n51_c;
                stage8_col111[1] = fa_s7_c111_n52_s;
                stage8_col112[0] = fa_s7_c111_n52_c;
                stage8_col112[1] = fa_s7_c112_n53_s;
                stage8_col113[0] = fa_s7_c112_n53_c;
                stage8_col113[1] = fa_s7_c113_n54_s;
                stage8_col114[0] = fa_s7_c113_n54_c;
                stage8_col114[1] = fa_s7_c114_n55_s;
                stage8_col115[0] = fa_s7_c114_n55_c;
                stage8_col115[1] = fa_s7_c115_n56_s;
                stage8_col116[0] = fa_s7_c115_n56_c;
                stage8_col116[1] = fa_s7_c116_n57_s;
                stage8_col117[0] = fa_s7_c116_n57_c;
                stage8_col117[1] = fa_s7_c117_n58_s;
                stage8_col118[0] = fa_s7_c117_n58_c;
                stage8_col118[1] = fa_s7_c118_n59_s;
                stage8_col119[0] = fa_s7_c118_n59_c;
                stage8_col119[1] = fa_s7_c119_n60_s;
                stage8_col120[0] = fa_s7_c119_n60_c;
                stage8_col120[1] = fa_s7_c120_n61_s;
                stage8_col121[0] = fa_s7_c120_n61_c;
                stage8_col121[1] = fa_s7_c121_n62_s;
                stage8_col122[0] = fa_s7_c121_n62_c;
                stage8_col122[1] = fa_s7_c122_n63_s;
                stage8_col123[0] = fa_s7_c122_n63_c;
                stage8_col123[1] = fa_s7_c123_n64_s;
                stage8_col124[0] = fa_s7_c123_n64_c;
                stage8_col124[1] = fa_s7_c124_n65_s;
                stage8_col125[0] = fa_s7_c124_n65_c;
                stage8_col125[1] = fa_s7_c125_n66_s;
                stage8_col126[0] = fa_s7_c125_n66_c;
                stage8_col126[1] = fa_s7_c126_n67_s;
                stage8_col127[0] = fa_s7_c126_n67_c;
                stage8_col127[1] = stage7_col127[0];
                stage8_col127[2] = stage7_col127[1];
                stage8_col127[3] = stage7_col127[2];
                stage8_col127[4] = stage7_col127[3];
                stage8_col127[5] = stage7_col127[4];
                stage8_col127[6] = stage7_col127[5];
                stage8_col127[7] = stage7_col127[6];
                stage8_col127[8] = stage7_col127[7];
                stage8_col127[9] = stage7_col127[8];
                stage8_col127[10] = stage7_col127[9];
                stage8_col127[11] = stage7_col127[10];
                stage8_col127[12] = stage7_col127[11];
                stage8_col127[13] = stage7_col127[12];
                stage8_col127[14] = stage7_col127[13];
                stage8_col127[15] = stage7_col127[14];
                stage8_col127[16] = stage7_col127[15];
                stage8_col127[17] = stage7_col127[16];
                stage8_col127[18] = stage7_col127[17];
                stage8_col127[19] = stage7_col127[18];
                stage8_col127[20] = stage7_col127[19];
                stage8_col127[21] = stage7_col127[20];
                stage8_col127[22] = stage7_col127[21];
                stage8_col127[23] = stage7_col127[22];
                stage8_col127[24] = stage7_col127[23];
                stage8_col127[25] = stage7_col127[24];
                stage8_col127[26] = stage7_col127[25];
                stage8_col127[27] = stage7_col127[26];
                stage8_col127[28] = stage7_col127[27];
                stage8_col127[29] = stage7_col127[28];
                stage8_col127[30] = stage7_col127[29];
                stage8_col127[31] = stage7_col127[30];
                stage8_col127[32] = stage7_col127[30];
                stage8_col127[33] = stage7_col127[30];
                stage8_col127[34] = stage7_col127[30];
                stage8_col127[35] = stage7_col127[30];
                stage8_col127[36] = stage7_col127[30];
                stage8_col127[37] = stage7_col127[30];
                stage8_col127[38] = stage7_col127[30];
                stage8_col127[39] = stage7_col127[30];
                stage8_col127[40] = stage7_col127[30];
                stage8_col127[41] = stage7_col127[30];
                stage8_col127[42] = stage7_col127[30];
                stage8_col127[43] = stage7_col127[30];
                stage8_col127[44] = stage7_col127[30];
                stage8_col127[45] = stage7_col127[30];
                stage8_col127[46] = stage7_col127[30];
                stage8_col127[47] = stage7_col127[30];
                stage8_col127[48] = stage7_col127[30];
                stage8_col127[49] = stage7_col127[30];
                stage8_col127[50] = stage7_col127[30];
                stage8_col127[51] = stage7_col127[30];
                stage8_col127[52] = stage7_col127[30];
                stage8_col127[53] = stage7_col127[30];
                stage8_col127[54] = stage7_col127[30];
                stage8_col127[55] = stage7_col127[30];
                stage8_col127[56] = stage7_col127[30];
                stage8_col127[57] = stage7_col127[30];
                stage8_col127[58] = stage7_col127[30];
                stage8_col127[59] = stage7_col127[30];
                stage8_col127[60] = stage7_col127[30];
                stage8_col127[61] = stage7_col127[30];
                stage8_col127[62] = stage7_col127[30];
            end
        end
    endgenerate

    // Final outputs (sum and carry)
    assign sum[0] = stage8_col0[0];
    assign carry[0] = 1'b0;
    assign sum[1] = stage8_col1[0];
    assign carry[1] = 1'b0;
    assign sum[2] = stage8_col2[0];
    assign carry[2] = 1'b0;
    assign sum[3] = stage8_col3[0];
    assign carry[3] = 1'b0;
    assign sum[4] = stage8_col4[0];
    assign carry[4] = 1'b0;
    assign sum[5] = stage8_col5[0];
    assign carry[5] = 1'b0;
    assign sum[6] = stage8_col6[0];
    assign carry[6] = 1'b0;
    assign sum[7] = stage8_col7[0];
    assign carry[7] = 1'b0;
    assign sum[8] = stage8_col8[0];
    assign carry[8] = stage8_col8[1];
    assign sum[9] = stage8_col9[0];
    assign carry[9] = 1'b0;
    assign sum[10] = stage8_col10[0];
    assign carry[10] = stage8_col10[1];
    assign sum[11] = stage8_col11[0];
    assign carry[11] = stage8_col11[1];
    assign sum[12] = stage8_col12[0];
    assign carry[12] = stage8_col12[1];
    assign sum[13] = stage8_col13[0];
    assign carry[13] = stage8_col13[1];
    assign sum[14] = stage8_col14[0];
    assign carry[14] = stage8_col14[1];
    assign sum[15] = stage8_col15[0];
    assign carry[15] = stage8_col15[1];
    assign sum[16] = stage8_col16[0];
    assign carry[16] = stage8_col16[1];
    assign sum[17] = stage8_col17[0];
    assign carry[17] = stage8_col17[1];
    assign sum[18] = stage8_col18[0];
    assign carry[18] = stage8_col18[1];
    assign sum[19] = stage8_col19[0];
    assign carry[19] = stage8_col19[1];
    assign sum[20] = stage8_col20[0];
    assign carry[20] = stage8_col20[1];
    assign sum[21] = stage8_col21[0];
    assign carry[21] = stage8_col21[1];
    assign sum[22] = stage8_col22[0];
    assign carry[22] = stage8_col22[1];
    assign sum[23] = stage8_col23[0];
    assign carry[23] = stage8_col23[1];
    assign sum[24] = stage8_col24[0];
    assign carry[24] = stage8_col24[1];
    assign sum[25] = stage8_col25[0];
    assign carry[25] = stage8_col25[1];
    assign sum[26] = stage8_col26[0];
    assign carry[26] = stage8_col26[1];
    assign sum[27] = stage8_col27[0];
    assign carry[27] = stage8_col27[1];
    assign sum[28] = stage8_col28[0];
    assign carry[28] = stage8_col28[1];
    assign sum[29] = stage8_col29[0];
    assign carry[29] = stage8_col29[1];
    assign sum[30] = stage8_col30[0];
    assign carry[30] = stage8_col30[1];
    assign sum[31] = stage8_col31[0];
    assign carry[31] = stage8_col31[1];
    assign sum[32] = stage8_col32[0];
    assign carry[32] = stage8_col32[1];
    assign sum[33] = stage8_col33[0];
    assign carry[33] = stage8_col33[1];
    assign sum[34] = stage8_col34[0];
    assign carry[34] = stage8_col34[1];
    assign sum[35] = stage8_col35[0];
    assign carry[35] = stage8_col35[1];
    assign sum[36] = stage8_col36[0];
    assign carry[36] = stage8_col36[1];
    assign sum[37] = stage8_col37[0];
    assign carry[37] = stage8_col37[1];
    assign sum[38] = stage8_col38[0];
    assign carry[38] = stage8_col38[1];
    assign sum[39] = stage8_col39[0];
    assign carry[39] = stage8_col39[1];
    assign sum[40] = stage8_col40[0];
    assign carry[40] = stage8_col40[1];
    assign sum[41] = stage8_col41[0];
    assign carry[41] = stage8_col41[1];
    assign sum[42] = stage8_col42[0];
    assign carry[42] = stage8_col42[1];
    assign sum[43] = stage8_col43[0];
    assign carry[43] = stage8_col43[1];
    assign sum[44] = stage8_col44[0];
    assign carry[44] = stage8_col44[1];
    assign sum[45] = stage8_col45[0];
    assign carry[45] = stage8_col45[1];
    assign sum[46] = stage8_col46[0];
    assign carry[46] = stage8_col46[1];
    assign sum[47] = stage8_col47[0];
    assign carry[47] = stage8_col47[1];
    assign sum[48] = stage8_col48[0];
    assign carry[48] = stage8_col48[1];
    assign sum[49] = stage8_col49[0];
    assign carry[49] = stage8_col49[1];
    assign sum[50] = stage8_col50[0];
    assign carry[50] = stage8_col50[1];
    assign sum[51] = stage8_col51[0];
    assign carry[51] = stage8_col51[1];
    assign sum[52] = stage8_col52[0];
    assign carry[52] = stage8_col52[1];
    assign sum[53] = stage8_col53[0];
    assign carry[53] = stage8_col53[1];
    assign sum[54] = stage8_col54[0];
    assign carry[54] = stage8_col54[1];
    assign sum[55] = stage8_col55[0];
    assign carry[55] = stage8_col55[1];
    assign sum[56] = stage8_col56[0];
    assign carry[56] = stage8_col56[1];
    assign sum[57] = stage8_col57[0];
    assign carry[57] = stage8_col57[1];
    assign sum[58] = stage8_col58[0];
    assign carry[58] = stage8_col58[1];
    assign sum[59] = stage8_col59[0];
    assign carry[59] = stage8_col59[1];
    assign sum[60] = stage8_col60[0];
    assign carry[60] = stage8_col60[1];
    assign sum[61] = stage8_col61[0];
    assign carry[61] = stage8_col61[1];
    assign sum[62] = stage8_col62[0];
    assign carry[62] = stage8_col62[1];
    assign sum[63] = stage8_col63[0];
    assign carry[63] = stage8_col63[1];
    assign sum[64] = stage8_col64[0];
    assign carry[64] = stage8_col64[1];
    assign sum[65] = stage8_col65[0];
    assign carry[65] = stage8_col65[1];
    assign sum[66] = stage8_col66[0];
    assign carry[66] = stage8_col66[1];
    assign sum[67] = stage8_col67[0];
    assign carry[67] = stage8_col67[1];
    assign sum[68] = stage8_col68[0];
    assign carry[68] = stage8_col68[1];
    assign sum[69] = stage8_col69[0];
    assign carry[69] = stage8_col69[1];
    assign sum[70] = stage8_col70[0];
    assign carry[70] = stage8_col70[1];
    assign sum[71] = stage8_col71[0];
    assign carry[71] = stage8_col71[1];
    assign sum[72] = stage8_col72[0];
    assign carry[72] = stage8_col72[1];
    assign sum[73] = stage8_col73[0];
    assign carry[73] = stage8_col73[1];
    assign sum[74] = stage8_col74[0];
    assign carry[74] = stage8_col74[1];
    assign sum[75] = stage8_col75[0];
    assign carry[75] = stage8_col75[1];
    assign sum[76] = stage8_col76[0];
    assign carry[76] = stage8_col76[1];
    assign sum[77] = stage8_col77[0];
    assign carry[77] = stage8_col77[1];
    assign sum[78] = stage8_col78[0];
    assign carry[78] = stage8_col78[1];
    assign sum[79] = stage8_col79[0];
    assign carry[79] = stage8_col79[1];
    assign sum[80] = stage8_col80[0];
    assign carry[80] = stage8_col80[1];
    assign sum[81] = stage8_col81[0];
    assign carry[81] = stage8_col81[1];
    assign sum[82] = stage8_col82[0];
    assign carry[82] = stage8_col82[1];
    assign sum[83] = stage8_col83[0];
    assign carry[83] = stage8_col83[1];
    assign sum[84] = stage8_col84[0];
    assign carry[84] = stage8_col84[1];
    assign sum[85] = stage8_col85[0];
    assign carry[85] = stage8_col85[1];
    assign sum[86] = stage8_col86[0];
    assign carry[86] = stage8_col86[1];
    assign sum[87] = stage8_col87[0];
    assign carry[87] = stage8_col87[1];
    assign sum[88] = stage8_col88[0];
    assign carry[88] = stage8_col88[1];
    assign sum[89] = stage8_col89[0];
    assign carry[89] = stage8_col89[1];
    assign sum[90] = stage8_col90[0];
    assign carry[90] = stage8_col90[1];
    assign sum[91] = stage8_col91[0];
    assign carry[91] = stage8_col91[1];
    assign sum[92] = stage8_col92[0];
    assign carry[92] = stage8_col92[1];
    assign sum[93] = stage8_col93[0];
    assign carry[93] = stage8_col93[1];
    assign sum[94] = stage8_col94[0];
    assign carry[94] = stage8_col94[1];
    assign sum[95] = stage8_col95[0];
    assign carry[95] = stage8_col95[1];
    assign sum[96] = stage8_col96[0];
    assign carry[96] = stage8_col96[1];
    assign sum[97] = stage8_col97[0];
    assign carry[97] = stage8_col97[1];
    assign sum[98] = stage8_col98[0];
    assign carry[98] = stage8_col98[1];
    assign sum[99] = stage8_col99[0];
    assign carry[99] = stage8_col99[1];
    assign sum[100] = stage8_col100[0];
    assign carry[100] = stage8_col100[1];
    assign sum[101] = stage8_col101[0];
    assign carry[101] = stage8_col101[1];
    assign sum[102] = stage8_col102[0];
    assign carry[102] = stage8_col102[1];
    assign sum[103] = stage8_col103[0];
    assign carry[103] = stage8_col103[1];
    assign sum[104] = stage8_col104[0];
    assign carry[104] = stage8_col104[1];
    assign sum[105] = stage8_col105[0];
    assign carry[105] = stage8_col105[1];
    assign sum[106] = stage8_col106[0];
    assign carry[106] = stage8_col106[1];
    assign sum[107] = stage8_col107[0];
    assign carry[107] = stage8_col107[1];
    assign sum[108] = stage8_col108[0];
    assign carry[108] = stage8_col108[1];
    assign sum[109] = stage8_col109[0];
    assign carry[109] = stage8_col109[1];
    assign sum[110] = stage8_col110[0];
    assign carry[110] = stage8_col110[1];
    assign sum[111] = stage8_col111[0];
    assign carry[111] = stage8_col111[1];
    assign sum[112] = stage8_col112[0];
    assign carry[112] = stage8_col112[1];
    assign sum[113] = stage8_col113[0];
    assign carry[113] = stage8_col113[1];
    assign sum[114] = stage8_col114[0];
    assign carry[114] = stage8_col114[1];
    assign sum[115] = stage8_col115[0];
    assign carry[115] = stage8_col115[1];
    assign sum[116] = stage8_col116[0];
    assign carry[116] = stage8_col116[1];
    assign sum[117] = stage8_col117[0];
    assign carry[117] = stage8_col117[1];
    assign sum[118] = stage8_col118[0];
    assign carry[118] = stage8_col118[1];
    assign sum[119] = stage8_col119[0];
    assign carry[119] = stage8_col119[1];
    assign sum[120] = stage8_col120[0];
    assign carry[120] = stage8_col120[1];
    assign sum[121] = stage8_col121[0];
    assign carry[121] = stage8_col121[1];
    assign sum[122] = stage8_col122[0];
    assign carry[122] = stage8_col122[1];
    assign sum[123] = stage8_col123[0];
    assign carry[123] = stage8_col123[1];
    assign sum[124] = stage8_col124[0];
    assign carry[124] = stage8_col124[1];
    assign sum[125] = stage8_col125[0];
    assign carry[125] = stage8_col125[1];
    assign sum[126] = stage8_col126[0];
    assign carry[126] = stage8_col126[1];
    // ERROR: More than 2 bits in final stage column 127
    assign sum[127] = ^(stage8_col127);
    assign carry[127] = 1'b0;

endmodule